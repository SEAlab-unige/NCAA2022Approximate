------------------------------------------------------------
-- Deeds (Digital Electronics Education and Design Suite)
-- VHDL Code generated on (4/30/2021, 4:28:02 PM)
--      by Deeds (Digital Circuit Simulator)(Deeds-DcS)
--      Ver. 2.40.330 (Jan 07, 2021)
-- Copyright (c) 2002-2020 University of Genoa, Italy
--      Web Site:  https://www.digitalelectronicsdeeds.com
------------------------------------------------------------

--------------------------------------------------------------------
LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY ROM256x16C200 IS         -- (programmable) ROM 256 x 16
  PORT( CS  : IN  std_logic;
        A00 : IN  std_logic;   -- ADR 7..0 (256 locations)
        A01 : IN  std_logic;
        A02 : IN  std_logic;
        A03 : IN  std_logic;
        A04 : IN  std_logic;
        A05 : IN  std_logic;
        A06 : IN  std_logic;
        A07 : IN  std_logic;
        D00 : OUT std_logic;   -- Data Output 15..00 (16-bits)
        D01 : OUT std_logic;
        D02 : OUT std_logic;
        D03 : OUT std_logic;
        D04 : OUT std_logic;
        D05 : OUT std_logic;
        D06 : OUT std_logic;
        D07 : OUT std_logic;
        D08 : OUT std_logic;
        D09 : OUT std_logic;
        D10 : OUT std_logic;
        D11 : OUT std_logic;
        D12 : OUT std_logic;
        D13 : OUT std_logic;
        D14 : OUT std_logic;
        D15 : OUT std_logic );
END ROM256x16C200;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF ROM256x16C200 IS
  --
  type ROM_Array is array (0 to 255) of std_logic_vector(15 downto 0);
  SIGNAL A : std_logic_vector( 7 downto 0);
  SIGNAL D : std_logic_vector(15 downto 0);

  -- ROM Memory Array ----------------------------------------------
  constant ROM_Cells: ROM_Array:= (
		00000 => "0000000000000011",
		00001 => "0000000000001111",
		00002 => "1111111111111111",
		00003 => "1111111111111111",
		00004 => "1111111111111111",
		00005 => "1111111111111111",
		00006 => "1111111111111111",
		00007 => "1111111111111111",
		00008 => "1111111111111111",
		00009 => "0011111111111111",
		00010 => "1111111111111111",
		00011 => "1111111111111111",
		00012 => "1111111111111111",
		00013 => "1111111111111111",
		00014 => "1111111111111111",
		00015 => "1111111111111111",
		00016 => "1111111111111111",
		00017 => "1111111111111111",
		00018 => "1111111111111111",
		00019 => "1111111111111111",
		00020 => "1111111111111111",
		00021 => "1111111111111111",
		00022 => "1111111111111111",
		00023 => "1111111111111111",
		00024 => "1111111111111111",
		00025 => "1111111111111111",
		00026 => "1111111111111111",
		00027 => "1101111111111111",
		00028 => "1111111111111111",
		00029 => "1111111111111111",
		00030 => "1111111111111111",
		00031 => "1111111111111111",
		00032 => "1111111111111111",
		00033 => "1101111111111111",
		00034 => "1111111111111111",
		00035 => "1111111111111111",
		00036 => "1111111111111111",
		00037 => "1111111111111111",
		00038 => "1111111111111111",
		00039 => "1111111111111111",
		00040 => "1111111111111111",
		00041 => "1111111111111111",
		00042 => "1111111111111111",
		00043 => "1111111111111111",
		00044 => "1111111111111111",
		00045 => "1111111111111111",
		00046 => "1111111111111111",
		00047 => "1111111111111111",
		00048 => "1111111111111111",
		00049 => "1111111111111111",
		00050 => "1111111111111111",
		00051 => "1111111111111111",
		00052 => "1111111111111111",
		00053 => "1111111111111111",
		00054 => "1111111111111111",
		00055 => "1111111111111111",
		00056 => "1111111111111111",
		00057 => "1111111111111111",
		00058 => "1111111111111111",
		00059 => "1111111111111111",
		00060 => "1111111111111111",
		00061 => "1111111111111111",
		00062 => "1111111111111111",
		00063 => "1111111111111111",
		00064 => "1111111111111111",
		00065 => "1111111111111111",
		00066 => "1111111111111111",
		00067 => "1111111111111111",
		00068 => "1111111111111111",
		00069 => "1111111111111111",
		00070 => "1111111111111111",
		00071 => "1111111111111111",
		00072 => "1111111111111111",
		00073 => "1111111111111111",
		00074 => "1111111111111111",
		00075 => "1111111111111111",
		00076 => "1111111111111111",
		00077 => "1111111111111111",
		00078 => "1111111111111111",
		00079 => "1111111111111111",
		00080 => "1111111111111111",
		00081 => "1111111111111111",
		00082 => "1111111111111111",
		00083 => "1111111111111111",
		00084 => "1111111111111111",
		00085 => "1111111111111111",
		00086 => "1111111111111111",
		00087 => "1111111111111111",
		00088 => "1111111111111111",
		00089 => "1111111111111111",
		00090 => "1111111111111111",
		00091 => "1111111111111111",
		00092 => "1111111111111111",
		00093 => "1111111111111111",
		00094 => "1111111111111111",
		00095 => "1111111111111111",
		00096 => "1111111111111111",
		00097 => "1111111111111111",
		00098 => "1111111111111111",
		00099 => "1111111111111111",
		00100 => "1111111111111111",
		00101 => "1111111111111111",
		00102 => "1111111111111111",
		00103 => "1111111111111111",
		00104 => "1111111111111111",
		00105 => "1111111111111111",
		00106 => "1111111111111111",
		00107 => "1111111111111111",
		00108 => "1111111111111111",
		00109 => "1111111111111111",
		00110 => "1111111111111111",
		00111 => "1111111111111111",
		00112 => "1111111111111111",
		00113 => "1111111111111111",
		00114 => "1111111111111111",
		00115 => "1111111111111111",
		00116 => "1111111111111111",
		00117 => "1111111111111111",
		00118 => "1111111111111111",
		00119 => "1111111111111111",
		00120 => "1111111111111111",
		00121 => "1111111111111111",
		00122 => "1111111111111111",
		00123 => "1111111111111111",
		00124 => "1111111111111111",
		00125 => "1111111111111111",
		00126 => "1111111111111111",
		00127 => "1111111111111111",
		00128 => "1111111111111111",
		00129 => "1111111111111111",
		00130 => "1111111111111111",
		00131 => "1111111111111111",
		00132 => "1111111111111111",
		00133 => "1111111111111111",
		00134 => "1111111111111111",
		00135 => "1111111111111111",
		00136 => "1111111111111111",
		00137 => "1111111111111111",
		00138 => "1111111111111111",
		00139 => "1111111111111111",
		00140 => "1111111111111111",
		00141 => "1111111111111111",
		00142 => "1111111111111111",
		00143 => "1111111111111111",
		00144 => "1111111111111111",
		00145 => "1111111111111111",
		00146 => "1111111111111111",
		00147 => "1111111111111111",
		00148 => "1111111111111111",
		00149 => "1111111111111111",
		00150 => "1111111111111111",
		00151 => "1111111111111111",
		00152 => "1111111111111111",
		00153 => "1111111111111111",
		00154 => "1111111111111111",
		00155 => "1111111111111111",
		00156 => "1111111111111111",
		00157 => "1111111111111111",
		00158 => "1111111111111111",
		00159 => "1111111111111111",
		00160 => "1111111111111111",
		00161 => "1111111111111111",
		00162 => "1111111111111111",
		00163 => "1111111111111111",
		00164 => "1111111111111111",
		00165 => "1111111111111111",
		00166 => "1111111111111111",
		00167 => "1111111111111111",
		00168 => "1111111111111111",
		00169 => "1111111111111111",
		00170 => "1111111111111111",
		00171 => "1111111111111111",
		00172 => "1111111111111111",
		00173 => "1111111111111111",
		00174 => "1111111111111111",
		00175 => "1111111111111111",
		00176 => "1111111111111111",
		00177 => "1111111111111111",
		00178 => "1111111111111111",
		00179 => "1111111111111111",
		00180 => "1111111111111111",
		00181 => "1111111111111111",
		00182 => "1111111111111111",
		00183 => "1111111111111111",
		00184 => "1111111111111111",
		00185 => "1111111111111111",
		00186 => "1111111111111111",
		00187 => "1111111111111111",
		00188 => "1111111111111111",
		00189 => "1111111111111111",
		00190 => "1111111111111111",
		00191 => "1111111111111111",
		00192 => "1111111111111111",
		00193 => "1111111111111111",
		00194 => "1111111111111111",
		00195 => "1111111111111111",
		00196 => "1111111111111111",
		00197 => "1111111111111111",
		00198 => "1111111111111111",
		00199 => "1111111111111111",
		00200 => "1111111111111111",
		00201 => "1111111111111111",
		00202 => "1111111111111111",
		00203 => "1111111111111111",
		00204 => "1111111111111111",
		00205 => "1111111111111111",
		00206 => "1111111111111111",
		00207 => "1111111111111111",
		00208 => "1111111111111111",
		00209 => "1111111111111111",
		00210 => "1111111111111111",
		00211 => "1111111111111111",
		00212 => "1111111111111111",
		00213 => "1111111111111111",
		00214 => "1111111111111111",
		00215 => "1111111111111111",
		00216 => "1111111111111111",
		00217 => "1111111111111111",
		00218 => "1111111111111111",
		00219 => "1111111111111111",
		00220 => "1111111111111111",
		00221 => "1111111111111111",
		00222 => "1111111111111111",
		00223 => "1111111111111111",
		00224 => "1111111111111111",
		00225 => "1111111111111111",
		00226 => "1111111111111111",
		00227 => "1111111111111111",
		00228 => "1111111111111111",
		00229 => "1111111111111111",
		00230 => "1111111111111111",
		00231 => "1111111111111111",
		00232 => "1111111111111111",
		00233 => "1111111111111111",
		00234 => "1111111111111111",
		00235 => "1111111111111111",
		00236 => "1111111111111111",
		00237 => "1111111111111111",
		00238 => "1111111111111111",
		00239 => "1111111111111111",
		00240 => "1111111111111111",
		00241 => "1111111111111111",
		00242 => "1111111111111111",
		00243 => "1111111111111111",
		00244 => "1111111111111111",
		00245 => "1111111111111111",
		00246 => "1111111111111111",
		00247 => "1111111111111111",
		00248 => "1111111111111111",
		00249 => "1111111111111111",
		00250 => "1111111111111111",
		00251 => "1111111111111111",
		00252 => "1111111111111111",
		00253 => "1111111111111111",
		00254 => "0000000000000000",
		00255 => "0000000000000000",
		OTHERS=> "1111111111111111"
		);

BEGIN
  A <= (A07 & A06 & A05 & A04 & A03 & A02 & A01 & A00);
  --
  PROCESS( CS, A )
  BEGIN
    if (CS = '1') then
          D <= ROM_Cells(to_integer(unsigned(A))); -- READ condition
    else  D <= (others => '0');                    -- Chip Select Off
    end if;
  END PROCESS;
  --
  D15 <= D(15); D14 <= D(14); D13 <= D(13); D12 <= D(12);
  D11 <= D(11); D10 <= D(10); D09 <= D(09); D08 <= D(08);
  D07 <= D(7);  D06 <= D(6);  D05 <= D(5);  D04 <= D(4);
  D03 <= D(3);  D02 <= D(2);  D01 <= D(1);  D00 <= D(0);
END behavioral;

--------------------------------------------------------------------
LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY ROM4kx8C1068 IS           -- (programmable) ROM 4k x 8
  PORT( CS  : IN  std_logic;
        A00 : IN  std_logic;   -- ADR 11..00 (4k locations)
        A01 : IN  std_logic;
        A02 : IN  std_logic;
        A03 : IN  std_logic;
        A04 : IN  std_logic;
        A05 : IN  std_logic;
        A06 : IN  std_logic;
        A07 : IN  std_logic;
        A08 : IN  std_logic;
        A09 : IN  std_logic;
        A10 : IN  std_logic;
        A11 : IN  std_logic;
        D00 : OUT std_logic;   -- Data Output 7..0 (8-bits)
        D01 : OUT std_logic;
        D02 : OUT std_logic;
        D03 : OUT std_logic;
        D04 : OUT std_logic;
        D05 : OUT std_logic;
        D06 : OUT std_logic;
        D07 : OUT std_logic );
END ROM4kx8C1068;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF ROM4kx8C1068 IS
  --
  type ROM_Array is array (0 to 4095) of std_logic_vector(7 downto 0);
  SIGNAL A : std_logic_vector(11 downto 0);
  SIGNAL D : std_logic_vector( 7 downto 0);

  -- ROM Memory Array ----------------------------------------------
  constant ROM_Cells: ROM_Array:= (
		00000 => "00000001",
		00001 => "00000010",
		00002 => "00000011",
		00003 => "00000100",
		00004 => "00000101",
		00005 => "00000110",
		00006 => "11111111",
		00007 => "11111111",
		00008 => "11111111",
		00009 => "11111111",
		00010 => "11111111",
		00011 => "11111111",
		00012 => "11111111",
		00013 => "11111111",
		00014 => "11111111",
		00015 => "11111111",
		00016 => "11111111",
		00017 => "11111111",
		00018 => "11111111",
		00019 => "11111111",
		00020 => "11111111",
		00021 => "11111111",
		00022 => "11111111",
		00023 => "11111111",
		00024 => "11111111",
		00025 => "11111111",
		00026 => "11111111",
		00027 => "11111111",
		00028 => "11111111",
		00029 => "11111111",
		00030 => "11111111",
		00031 => "11111111",
		00032 => "11111111",
		00033 => "11111111",
		00034 => "11111111",
		00035 => "11111111",
		00036 => "11111111",
		00037 => "11111111",
		00038 => "11111111",
		00039 => "11111111",
		00040 => "11111111",
		00041 => "11111111",
		00042 => "11111111",
		00043 => "11111111",
		00044 => "11111111",
		00045 => "11111111",
		00046 => "11111111",
		00047 => "11111111",
		00048 => "11111111",
		00049 => "11111111",
		00050 => "11111111",
		00051 => "11111111",
		00052 => "11111111",
		00053 => "11111111",
		00054 => "11111111",
		00055 => "11111111",
		00056 => "11111111",
		00057 => "11111111",
		00058 => "11111111",
		00059 => "11111111",
		00060 => "11111111",
		00061 => "11111111",
		00062 => "11111111",
		00063 => "11111111",
		00064 => "11111111",
		00065 => "11111111",
		00066 => "11111111",
		00067 => "11111111",
		00068 => "11111111",
		00069 => "11111111",
		00070 => "11111111",
		00071 => "11111111",
		00072 => "11111111",
		00073 => "11111111",
		00074 => "11111111",
		00075 => "11111111",
		00076 => "11111111",
		00077 => "11111111",
		00078 => "11111111",
		00079 => "11111111",
		00080 => "11111111",
		00081 => "11111111",
		00082 => "11111111",
		00083 => "11111111",
		00084 => "11111111",
		00085 => "11111111",
		00086 => "11111111",
		00087 => "11111111",
		00088 => "11111111",
		00089 => "11111111",
		00090 => "11111111",
		00091 => "11111111",
		00092 => "11111111",
		00093 => "11111111",
		00094 => "11111111",
		00095 => "11111111",
		00096 => "11111111",
		00097 => "11111111",
		00098 => "11111111",
		00099 => "11111111",
		00100 => "11111111",
		00101 => "11111111",
		00102 => "11111111",
		00103 => "11111111",
		00104 => "11111111",
		00105 => "11111111",
		00106 => "11111111",
		00107 => "11111111",
		00108 => "11111111",
		00109 => "11111111",
		00110 => "11111111",
		00111 => "11111111",
		00112 => "11111111",
		00113 => "11111111",
		00114 => "11111111",
		00115 => "11111111",
		00116 => "11111111",
		00117 => "11111111",
		00118 => "11111111",
		00119 => "11111111",
		00120 => "11111111",
		00121 => "11111111",
		00122 => "11111111",
		00123 => "11111111",
		00124 => "11111111",
		00125 => "11111111",
		00126 => "11111111",
		00127 => "11111111",
		00128 => "11111111",
		00129 => "11111111",
		00130 => "11111111",
		00131 => "11111111",
		00132 => "11111111",
		00133 => "11111111",
		00134 => "11111111",
		00135 => "11111111",
		00136 => "11111111",
		00137 => "11111111",
		00138 => "11111111",
		00139 => "11111111",
		00140 => "11111111",
		00141 => "11111111",
		00142 => "11111111",
		00143 => "11111111",
		00144 => "11111111",
		00145 => "11111111",
		00146 => "11111111",
		00147 => "11111111",
		00148 => "11111111",
		00149 => "11111111",
		00150 => "11111111",
		00151 => "11111111",
		00152 => "11111111",
		00153 => "11111111",
		00154 => "11111111",
		00155 => "11111111",
		00156 => "11111111",
		00157 => "11111111",
		00158 => "11111111",
		00159 => "11111111",
		00160 => "11111111",
		00161 => "11111111",
		00162 => "11111111",
		00163 => "11111111",
		00164 => "11111111",
		00165 => "11111111",
		00166 => "11111111",
		00167 => "11111111",
		00168 => "11111111",
		00169 => "11111111",
		00170 => "11111111",
		00171 => "11111111",
		00172 => "11111111",
		00173 => "11111111",
		00174 => "11111111",
		00175 => "11111111",
		00176 => "11111111",
		00177 => "11111111",
		00178 => "11111111",
		00179 => "11111111",
		00180 => "11111111",
		00181 => "11111111",
		00182 => "11111111",
		00183 => "11111111",
		00184 => "11111111",
		00185 => "11111111",
		00186 => "11111111",
		00187 => "11111111",
		00188 => "11111111",
		00189 => "11111111",
		00190 => "11111111",
		00191 => "11111111",
		00192 => "11111111",
		00193 => "11111111",
		00194 => "11111111",
		00195 => "11111111",
		00196 => "11111111",
		00197 => "11111111",
		00198 => "11111111",
		00199 => "11111111",
		00200 => "11111111",
		00201 => "11111111",
		00202 => "11111111",
		00203 => "11111111",
		00204 => "11111111",
		00205 => "11111111",
		00206 => "11111111",
		00207 => "11111111",
		00208 => "11111111",
		00209 => "11111111",
		00210 => "11111111",
		00211 => "11111111",
		00212 => "11111111",
		00213 => "11111111",
		00214 => "11111111",
		00215 => "11111111",
		00216 => "11111111",
		00217 => "11111111",
		00218 => "11111111",
		00219 => "11111111",
		00220 => "11111111",
		00221 => "11111111",
		00222 => "11111111",
		00223 => "11111111",
		00224 => "11111111",
		00225 => "11111111",
		00226 => "11111111",
		00227 => "11111111",
		00228 => "11111111",
		00229 => "11111111",
		00230 => "11111111",
		00231 => "11111111",
		00232 => "11111111",
		00233 => "11111111",
		00234 => "11111111",
		00235 => "11111111",
		00236 => "11111111",
		00237 => "11111111",
		00238 => "11111111",
		00239 => "11111111",
		00240 => "11111111",
		00241 => "11111111",
		00242 => "11111111",
		00243 => "11111111",
		00244 => "11111111",
		00245 => "11111111",
		00246 => "11111111",
		00247 => "11111111",
		00248 => "11111111",
		00249 => "11111111",
		00250 => "11111111",
		00251 => "11111111",
		00252 => "11111111",
		00253 => "11111111",
		00254 => "11111111",
		00255 => "11111111",
		00256 => "11111111",
		00257 => "11111111",
		00258 => "11111111",
		00259 => "11111111",
		00260 => "11111111",
		00261 => "11111111",
		00262 => "11111111",
		00263 => "11111111",
		00264 => "11111111",
		00265 => "11111111",
		00266 => "11111111",
		00267 => "11111111",
		00268 => "11111111",
		00269 => "11111111",
		00270 => "11111111",
		00271 => "11111111",
		00272 => "11111111",
		00273 => "11111111",
		00274 => "11111111",
		00275 => "11111111",
		00276 => "11111111",
		00277 => "11111111",
		00278 => "11111111",
		00279 => "11111111",
		00280 => "11111111",
		00281 => "11111111",
		00282 => "11111111",
		00283 => "11111111",
		00284 => "11111111",
		00285 => "11111111",
		00286 => "11111111",
		00287 => "11111111",
		00288 => "11111111",
		00289 => "11111111",
		00290 => "11111111",
		00291 => "11111111",
		00292 => "11111111",
		00293 => "11111111",
		00294 => "11111111",
		00295 => "11111111",
		00296 => "11111111",
		00297 => "11111111",
		00298 => "11111111",
		00299 => "11111111",
		00300 => "11111111",
		00301 => "11111111",
		00302 => "11111111",
		00303 => "11111111",
		00304 => "11111111",
		00305 => "11111111",
		00306 => "11111111",
		00307 => "11111111",
		00308 => "11111111",
		00309 => "11111111",
		00310 => "11111111",
		00311 => "11111111",
		00312 => "11111111",
		00313 => "11111111",
		00314 => "11111111",
		00315 => "11111111",
		00316 => "11111111",
		00317 => "11111111",
		00318 => "11111111",
		00319 => "11111111",
		00320 => "11111111",
		00321 => "11111111",
		00322 => "11111111",
		00323 => "11111111",
		00324 => "11111111",
		00325 => "11111111",
		00326 => "11111111",
		00327 => "11111111",
		00328 => "11111111",
		00329 => "11111111",
		00330 => "11111111",
		00331 => "11111111",
		00332 => "11111111",
		00333 => "11111111",
		00334 => "11111111",
		00335 => "11111111",
		00336 => "11111111",
		00337 => "11111111",
		00338 => "11111111",
		00339 => "11111111",
		00340 => "11111111",
		00341 => "11111111",
		00342 => "11111111",
		00343 => "11111111",
		00344 => "11111111",
		00345 => "11111111",
		00346 => "11111111",
		00347 => "11111111",
		00348 => "11111111",
		00349 => "11111111",
		00350 => "11111111",
		00351 => "11111111",
		00352 => "11111111",
		00353 => "11111111",
		00354 => "11111111",
		00355 => "11111111",
		00356 => "11111111",
		00357 => "11111111",
		00358 => "11111111",
		00359 => "11111111",
		00360 => "11111111",
		00361 => "11111111",
		00362 => "11111111",
		00363 => "11111111",
		00364 => "11111111",
		00365 => "11111111",
		00366 => "11111111",
		00367 => "11111111",
		00368 => "11111111",
		00369 => "11111111",
		00370 => "11111111",
		00371 => "11111111",
		00372 => "11111111",
		00373 => "11111111",
		00374 => "11111111",
		00375 => "11111111",
		00376 => "11111111",
		00377 => "11111111",
		00378 => "11111111",
		00379 => "11111111",
		00380 => "11111111",
		00381 => "11111111",
		00382 => "11111111",
		00383 => "11111111",
		00384 => "11111111",
		00385 => "11111111",
		00386 => "11111111",
		00387 => "11111111",
		00388 => "11111111",
		00389 => "11111111",
		00390 => "11111111",
		00391 => "11111111",
		00392 => "11111111",
		00393 => "11111111",
		00394 => "11111111",
		00395 => "11111111",
		00396 => "11111111",
		00397 => "11111111",
		00398 => "11111111",
		00399 => "11111111",
		00400 => "11111111",
		00401 => "11111111",
		00402 => "11111111",
		00403 => "11111111",
		00404 => "11111111",
		00405 => "11111111",
		00406 => "11111111",
		00407 => "11111111",
		00408 => "11111111",
		00409 => "11111111",
		00410 => "11111111",
		00411 => "11111111",
		00412 => "11111111",
		00413 => "11111111",
		00414 => "11111111",
		00415 => "11111111",
		00416 => "11111111",
		00417 => "11111111",
		00418 => "11111111",
		00419 => "11111111",
		00420 => "11111111",
		00421 => "11111111",
		00422 => "11111111",
		00423 => "11111111",
		00424 => "11111111",
		00425 => "11111111",
		00426 => "11111111",
		00427 => "11111111",
		00428 => "11111111",
		00429 => "11111111",
		00430 => "11111111",
		00431 => "11111111",
		00432 => "11111111",
		00433 => "11111111",
		00434 => "11111111",
		00435 => "11111111",
		00436 => "11111111",
		00437 => "11111111",
		00438 => "11111111",
		00439 => "11111111",
		00440 => "11111111",
		00441 => "11111111",
		00442 => "11111111",
		00443 => "11111111",
		00444 => "11111111",
		00445 => "11111111",
		00446 => "11111111",
		00447 => "11111111",
		00448 => "11111111",
		00449 => "11111111",
		00450 => "11111111",
		00451 => "11111111",
		00452 => "11111111",
		00453 => "11111111",
		00454 => "11111111",
		00455 => "11111111",
		00456 => "11111111",
		00457 => "11111111",
		00458 => "11111111",
		00459 => "11111111",
		00460 => "11111111",
		00461 => "11111111",
		00462 => "11111111",
		00463 => "11111111",
		00464 => "11111111",
		00465 => "11111111",
		00466 => "11111111",
		00467 => "11111111",
		00468 => "11111111",
		00469 => "11111111",
		00470 => "11111111",
		00471 => "11111111",
		00472 => "11111111",
		00473 => "11111111",
		00474 => "11111111",
		00475 => "11111111",
		00476 => "11111111",
		00477 => "11111111",
		00478 => "11111111",
		00479 => "11111111",
		00480 => "11111111",
		00481 => "11111111",
		00482 => "11111111",
		00483 => "11111111",
		00484 => "11111111",
		00485 => "11111111",
		00486 => "11111111",
		00487 => "11111111",
		00488 => "11111111",
		00489 => "11111111",
		00490 => "11111111",
		00491 => "11111111",
		00492 => "11111111",
		00493 => "11111111",
		00494 => "11111111",
		00495 => "11111111",
		00496 => "11111111",
		00497 => "11111111",
		00498 => "11111111",
		00499 => "11111111",
		00500 => "11111111",
		00501 => "11111111",
		00502 => "11111111",
		00503 => "11111111",
		00504 => "11111111",
		00505 => "11111111",
		00506 => "11111111",
		00507 => "11111111",
		00508 => "11111111",
		00509 => "11111111",
		00510 => "11111111",
		00511 => "11111111",
		00512 => "11111111",
		00513 => "11111111",
		00514 => "11111111",
		00515 => "11111111",
		00516 => "11111111",
		00517 => "11111111",
		00518 => "11111111",
		00519 => "11111111",
		00520 => "11111111",
		00521 => "11111111",
		00522 => "11111111",
		00523 => "11111111",
		00524 => "11111111",
		00525 => "11111111",
		00526 => "11111111",
		00527 => "11111111",
		00528 => "11111111",
		00529 => "11111111",
		00530 => "11111111",
		00531 => "11111111",
		00532 => "11111111",
		00533 => "11111111",
		00534 => "11111111",
		00535 => "11111111",
		00536 => "11111111",
		00537 => "11111111",
		00538 => "11111111",
		00539 => "11111111",
		00540 => "11111111",
		00541 => "11111111",
		00542 => "11111111",
		00543 => "11111111",
		00544 => "11111111",
		00545 => "11111111",
		00546 => "11111111",
		00547 => "11111111",
		00548 => "11111111",
		00549 => "11111111",
		00550 => "11111111",
		00551 => "11111111",
		00552 => "11111111",
		00553 => "11111111",
		00554 => "11111111",
		00555 => "11111111",
		00556 => "11111111",
		00557 => "11111111",
		00558 => "11111111",
		00559 => "11111111",
		00560 => "11111111",
		00561 => "11111111",
		00562 => "11111111",
		00563 => "11111111",
		00564 => "11111111",
		00565 => "11111111",
		00566 => "11111111",
		00567 => "11111111",
		00568 => "11111111",
		00569 => "11111111",
		00570 => "11111111",
		00571 => "11111111",
		00572 => "11111111",
		00573 => "11111111",
		00574 => "11111111",
		00575 => "11111111",
		00576 => "11111111",
		00577 => "11111111",
		00578 => "11111111",
		00579 => "11111111",
		00580 => "11111111",
		00581 => "11111111",
		00582 => "11111111",
		00583 => "11111111",
		00584 => "11111111",
		00585 => "11111111",
		00586 => "11111111",
		00587 => "11111111",
		00588 => "11111111",
		00589 => "11111111",
		00590 => "11111111",
		00591 => "11111111",
		00592 => "11111111",
		00593 => "11111111",
		00594 => "11111111",
		00595 => "11111111",
		00596 => "11111111",
		00597 => "11111111",
		00598 => "11111111",
		00599 => "11111111",
		00600 => "11111111",
		00601 => "11111111",
		00602 => "11111111",
		00603 => "11111111",
		00604 => "11111111",
		00605 => "11111111",
		00606 => "11111111",
		00607 => "11111111",
		00608 => "11111111",
		00609 => "11111111",
		00610 => "11111111",
		00611 => "11111111",
		00612 => "11111111",
		00613 => "11111111",
		00614 => "11111111",
		00615 => "11111111",
		00616 => "11111111",
		00617 => "11111111",
		00618 => "11111111",
		00619 => "11111111",
		00620 => "11111111",
		00621 => "11111111",
		00622 => "11111111",
		00623 => "11111111",
		00624 => "11111111",
		00625 => "11111111",
		00626 => "11111111",
		00627 => "11111111",
		00628 => "11111111",
		00629 => "11111111",
		00630 => "11111111",
		00631 => "11111111",
		00632 => "11111111",
		00633 => "11111111",
		00634 => "11111111",
		00635 => "11111111",
		00636 => "11111111",
		00637 => "11111111",
		00638 => "11111111",
		00639 => "11111111",
		00640 => "11111111",
		00641 => "11111111",
		00642 => "11111111",
		00643 => "11111111",
		00644 => "11111111",
		00645 => "11111111",
		00646 => "11111111",
		00647 => "11111111",
		00648 => "11111111",
		00649 => "11111111",
		00650 => "11111111",
		00651 => "11111111",
		00652 => "11111111",
		00653 => "11111111",
		00654 => "11111111",
		00655 => "11111111",
		00656 => "11111111",
		00657 => "11111111",
		00658 => "11111111",
		00659 => "11111111",
		00660 => "11111111",
		00661 => "11111111",
		00662 => "11111111",
		00663 => "11111111",
		00664 => "11111111",
		00665 => "11111111",
		00666 => "11111111",
		00667 => "11111111",
		00668 => "11111111",
		00669 => "11111111",
		00670 => "11111111",
		00671 => "11111111",
		00672 => "11111111",
		00673 => "11111111",
		00674 => "11111111",
		00675 => "11111111",
		00676 => "11111111",
		00677 => "11111111",
		00678 => "11111111",
		00679 => "11111111",
		00680 => "11111111",
		00681 => "11111111",
		00682 => "11111111",
		00683 => "11111111",
		00684 => "11111111",
		00685 => "11111111",
		00686 => "11111111",
		00687 => "11111111",
		00688 => "11111111",
		00689 => "11111111",
		00690 => "11111111",
		00691 => "11111111",
		00692 => "11111111",
		00693 => "11111111",
		00694 => "11111111",
		00695 => "11111111",
		00696 => "11111111",
		00697 => "11111111",
		00698 => "11111111",
		00699 => "11111111",
		00700 => "11111111",
		00701 => "11111111",
		00702 => "11111111",
		00703 => "11111111",
		00704 => "11111111",
		00705 => "11111111",
		00706 => "11111111",
		00707 => "11111111",
		00708 => "11111111",
		00709 => "11111111",
		00710 => "11111111",
		00711 => "11111111",
		00712 => "11111111",
		00713 => "11111111",
		00714 => "11111111",
		00715 => "11111111",
		00716 => "11111111",
		00717 => "11111111",
		00718 => "11111111",
		00719 => "11111111",
		00720 => "11111111",
		00721 => "11111111",
		00722 => "11111111",
		00723 => "11111111",
		00724 => "11111111",
		00725 => "11111111",
		00726 => "11111111",
		00727 => "11111111",
		00728 => "11111111",
		00729 => "11111111",
		00730 => "11111111",
		00731 => "11111111",
		00732 => "11111111",
		00733 => "11111111",
		00734 => "11111111",
		00735 => "11111111",
		00736 => "11111111",
		00737 => "11111111",
		00738 => "11111111",
		00739 => "11111111",
		00740 => "11111111",
		00741 => "11111111",
		00742 => "11111111",
		00743 => "11111111",
		00744 => "11111111",
		00745 => "11111111",
		00746 => "11111111",
		00747 => "11111111",
		00748 => "11111111",
		00749 => "11111111",
		00750 => "11111111",
		00751 => "11111111",
		00752 => "11111111",
		00753 => "11111111",
		00754 => "11111111",
		00755 => "11111111",
		00756 => "11111111",
		00757 => "11111111",
		00758 => "11111111",
		00759 => "11111111",
		00760 => "11111111",
		00761 => "11111111",
		00762 => "11111111",
		00763 => "11111111",
		00764 => "11111111",
		00765 => "11111111",
		00766 => "11111111",
		00767 => "11111111",
		00768 => "11111111",
		00769 => "11111111",
		00770 => "11111111",
		00771 => "11111111",
		00772 => "11111111",
		00773 => "11111111",
		00774 => "11111111",
		00775 => "11111111",
		00776 => "11111111",
		00777 => "11111111",
		00778 => "11111111",
		00779 => "11111111",
		00780 => "11111111",
		00781 => "11111111",
		00782 => "11111111",
		00783 => "11111111",
		00784 => "11111111",
		00785 => "11111111",
		00786 => "11111111",
		00787 => "11111111",
		00788 => "11111111",
		00789 => "11111111",
		00790 => "11111111",
		00791 => "11111111",
		00792 => "11111111",
		00793 => "11111111",
		00794 => "11111111",
		00795 => "11111111",
		00796 => "11111111",
		00797 => "11111111",
		00798 => "11111111",
		00799 => "11111111",
		00800 => "11111111",
		00801 => "11111111",
		00802 => "11111111",
		00803 => "11111111",
		00804 => "11111111",
		00805 => "11111111",
		00806 => "11111111",
		00807 => "11111111",
		00808 => "11111111",
		00809 => "11111111",
		00810 => "11111111",
		00811 => "11111111",
		00812 => "11111111",
		00813 => "11111111",
		00814 => "11111111",
		00815 => "11111111",
		00816 => "11111111",
		00817 => "11111111",
		00818 => "11111111",
		00819 => "11111111",
		00820 => "11111111",
		00821 => "11111111",
		00822 => "11111111",
		00823 => "11111111",
		00824 => "11111111",
		00825 => "11111111",
		00826 => "11111111",
		00827 => "11111111",
		00828 => "11111111",
		00829 => "11111111",
		00830 => "11111111",
		00831 => "11111111",
		00832 => "11111111",
		00833 => "11111111",
		00834 => "11111111",
		00835 => "11111111",
		00836 => "11111111",
		00837 => "11111111",
		00838 => "11111111",
		00839 => "11111111",
		00840 => "11111111",
		00841 => "11111111",
		00842 => "11111111",
		00843 => "11111111",
		00844 => "11111111",
		00845 => "11111111",
		00846 => "11111111",
		00847 => "11111111",
		00848 => "11111111",
		00849 => "11111111",
		00850 => "11111111",
		00851 => "11111111",
		00852 => "11111111",
		00853 => "11111111",
		00854 => "11111111",
		00855 => "11111111",
		00856 => "11111111",
		00857 => "11111111",
		00858 => "11111111",
		00859 => "11111111",
		00860 => "11111111",
		00861 => "11111111",
		00862 => "11111111",
		00863 => "11111111",
		00864 => "11111111",
		00865 => "11111111",
		00866 => "11111111",
		00867 => "11111111",
		00868 => "11111111",
		00869 => "11111111",
		00870 => "11111111",
		00871 => "11111111",
		00872 => "11111111",
		00873 => "11111111",
		00874 => "11111111",
		00875 => "11111111",
		00876 => "11111111",
		00877 => "11111111",
		00878 => "11111111",
		00879 => "11111111",
		00880 => "11111111",
		00881 => "11111111",
		00882 => "11111111",
		00883 => "11111111",
		00884 => "11111111",
		00885 => "11111111",
		00886 => "11111111",
		00887 => "11111111",
		00888 => "11111111",
		00889 => "11111111",
		00890 => "11111111",
		00891 => "11111111",
		00892 => "11111111",
		00893 => "11111111",
		00894 => "11111111",
		00895 => "11111111",
		00896 => "11111111",
		00897 => "11111111",
		00898 => "11111111",
		00899 => "11111111",
		00900 => "11111111",
		00901 => "11111111",
		00902 => "11111111",
		00903 => "11111111",
		00904 => "11111111",
		00905 => "11111111",
		00906 => "11111111",
		00907 => "11111111",
		00908 => "11111111",
		00909 => "11111111",
		00910 => "11111111",
		00911 => "11111111",
		00912 => "11111111",
		00913 => "11111111",
		00914 => "11111111",
		00915 => "11111111",
		00916 => "11111111",
		00917 => "11111111",
		00918 => "11111111",
		00919 => "11111111",
		00920 => "11111111",
		00921 => "11111111",
		00922 => "11111111",
		00923 => "11111111",
		00924 => "11111111",
		00925 => "11111111",
		00926 => "11111111",
		00927 => "11111111",
		00928 => "11111111",
		00929 => "11111111",
		00930 => "11111111",
		00931 => "11111111",
		00932 => "11111111",
		00933 => "11111111",
		00934 => "11111111",
		00935 => "11111111",
		00936 => "11111111",
		00937 => "11111111",
		00938 => "11111111",
		00939 => "11111111",
		00940 => "11111111",
		00941 => "11111111",
		00942 => "11111111",
		00943 => "11111111",
		00944 => "11111111",
		00945 => "11111111",
		00946 => "11111111",
		00947 => "11111111",
		00948 => "11111111",
		00949 => "11111111",
		00950 => "11111111",
		00951 => "11111111",
		00952 => "11111111",
		00953 => "11111111",
		00954 => "11111111",
		00955 => "11111111",
		00956 => "11111111",
		00957 => "11111111",
		00958 => "11111111",
		00959 => "11111111",
		00960 => "11111111",
		00961 => "11111111",
		00962 => "11111111",
		00963 => "11111111",
		00964 => "11111111",
		00965 => "11111111",
		00966 => "11111111",
		00967 => "11111111",
		00968 => "11111111",
		00969 => "11111111",
		00970 => "11111111",
		00971 => "11111111",
		00972 => "11111111",
		00973 => "11111111",
		00974 => "11111111",
		00975 => "11111111",
		00976 => "11111111",
		00977 => "11111111",
		00978 => "11111111",
		00979 => "11111111",
		00980 => "11111111",
		00981 => "11111111",
		00982 => "11111111",
		00983 => "11111111",
		00984 => "11111111",
		00985 => "11111111",
		00986 => "11111111",
		00987 => "11111111",
		00988 => "11111111",
		00989 => "11111111",
		00990 => "11111111",
		00991 => "11111111",
		00992 => "11111111",
		00993 => "11111111",
		00994 => "11111111",
		00995 => "11111111",
		00996 => "11111111",
		00997 => "11111111",
		00998 => "11111111",
		00999 => "11111111",
		01000 => "11111111",
		01001 => "11111111",
		01002 => "11111111",
		01003 => "11111111",
		01004 => "11111111",
		01005 => "11111111",
		01006 => "11111111",
		01007 => "11111111",
		01008 => "11111111",
		01009 => "11111111",
		01010 => "11111111",
		01011 => "11111111",
		01012 => "11111111",
		01013 => "11111111",
		01014 => "11111111",
		01015 => "11111111",
		01016 => "11111111",
		01017 => "11111111",
		01018 => "11111111",
		01019 => "11111111",
		01020 => "11111111",
		01021 => "11111111",
		01022 => "11111111",
		01023 => "11111111",
		01024 => "11111111",
		01025 => "11111111",
		01026 => "11111111",
		01027 => "11111111",
		01028 => "11111111",
		01029 => "11111111",
		01030 => "11111111",
		01031 => "11111111",
		01032 => "11111111",
		01033 => "11111111",
		01034 => "11111111",
		01035 => "11111111",
		01036 => "11111111",
		01037 => "11111111",
		01038 => "11111111",
		01039 => "11111111",
		01040 => "11111111",
		01041 => "11111111",
		01042 => "11111111",
		01043 => "11111111",
		01044 => "11111111",
		01045 => "11111111",
		01046 => "11111111",
		01047 => "11111111",
		01048 => "11111111",
		01049 => "11111111",
		01050 => "11111111",
		01051 => "11111111",
		01052 => "11111111",
		01053 => "11111111",
		01054 => "11111111",
		01055 => "11111111",
		01056 => "11111111",
		01057 => "11111111",
		01058 => "11111111",
		01059 => "11111111",
		01060 => "11111111",
		01061 => "11111111",
		01062 => "11111111",
		01063 => "11111111",
		01064 => "11111111",
		01065 => "11111111",
		01066 => "11111111",
		01067 => "11111111",
		01068 => "11111111",
		01069 => "11111111",
		01070 => "11111111",
		01071 => "11111111",
		01072 => "11111111",
		01073 => "11111111",
		01074 => "11111111",
		01075 => "11111111",
		01076 => "11111111",
		01077 => "11111111",
		01078 => "11111111",
		01079 => "11111111",
		01080 => "11111111",
		01081 => "11111111",
		01082 => "11111111",
		01083 => "11111111",
		01084 => "11111111",
		01085 => "11111111",
		01086 => "11111111",
		01087 => "11111111",
		01088 => "11111111",
		01089 => "11111111",
		01090 => "11111111",
		01091 => "11111111",
		01092 => "11111111",
		01093 => "11111111",
		01094 => "11111111",
		01095 => "11111111",
		01096 => "11111111",
		01097 => "11111111",
		01098 => "11111111",
		01099 => "11111111",
		01100 => "11111111",
		01101 => "11111111",
		01102 => "11111111",
		01103 => "11111111",
		01104 => "11111111",
		01105 => "11111111",
		01106 => "11111111",
		01107 => "11111111",
		01108 => "11111111",
		01109 => "11111111",
		01110 => "11111111",
		01111 => "11111111",
		01112 => "11111111",
		01113 => "11111111",
		01114 => "11111111",
		01115 => "11111111",
		01116 => "11111111",
		01117 => "11111111",
		01118 => "11111111",
		01119 => "11111111",
		01120 => "11111111",
		01121 => "11111111",
		01122 => "11111111",
		01123 => "11111111",
		01124 => "11111111",
		01125 => "11111111",
		01126 => "11111111",
		01127 => "11111111",
		01128 => "11111111",
		01129 => "11111111",
		01130 => "11111111",
		01131 => "11111111",
		01132 => "11111111",
		01133 => "11111111",
		01134 => "11111111",
		01135 => "11111111",
		01136 => "11111111",
		01137 => "11111111",
		01138 => "11111111",
		01139 => "11111111",
		01140 => "11111111",
		01141 => "11111111",
		01142 => "11111111",
		01143 => "11111111",
		01144 => "11111111",
		01145 => "11111111",
		01146 => "11111111",
		01147 => "11111111",
		01148 => "11111111",
		01149 => "11111111",
		01150 => "11111111",
		01151 => "11111111",
		01152 => "11111111",
		01153 => "11111111",
		01154 => "11111111",
		01155 => "11111111",
		01156 => "11111111",
		01157 => "11111111",
		01158 => "11111111",
		01159 => "11111111",
		01160 => "11111111",
		01161 => "11111111",
		01162 => "11111111",
		01163 => "11111111",
		01164 => "11111111",
		01165 => "11111111",
		01166 => "11111111",
		01167 => "11111111",
		01168 => "11111111",
		01169 => "11111111",
		01170 => "11111111",
		01171 => "11111111",
		01172 => "11111111",
		01173 => "11111111",
		01174 => "11111111",
		01175 => "11111111",
		01176 => "11111111",
		01177 => "11111111",
		01178 => "11111111",
		01179 => "11111111",
		01180 => "11111111",
		01181 => "11111111",
		01182 => "11111111",
		01183 => "11111111",
		01184 => "11111111",
		01185 => "11111111",
		01186 => "11111111",
		01187 => "11111111",
		01188 => "11111111",
		01189 => "11111111",
		01190 => "11111111",
		01191 => "11111111",
		01192 => "11111111",
		01193 => "11111111",
		01194 => "11111111",
		01195 => "11111111",
		01196 => "11111111",
		01197 => "11111111",
		01198 => "11111111",
		01199 => "11111111",
		01200 => "11111111",
		01201 => "11111111",
		01202 => "11111111",
		01203 => "11111111",
		01204 => "11111111",
		01205 => "11111111",
		01206 => "11111111",
		01207 => "11111111",
		01208 => "11111111",
		01209 => "11111111",
		01210 => "11111111",
		01211 => "11111111",
		01212 => "11111111",
		01213 => "11111111",
		01214 => "11111111",
		01215 => "11111111",
		01216 => "11111111",
		01217 => "11111111",
		01218 => "11111111",
		01219 => "11111111",
		01220 => "11111111",
		01221 => "11111111",
		01222 => "11111111",
		01223 => "11111111",
		01224 => "11111111",
		01225 => "11111111",
		01226 => "11111111",
		01227 => "11111111",
		01228 => "11111111",
		01229 => "11111111",
		01230 => "11111111",
		01231 => "11111111",
		01232 => "11111111",
		01233 => "11111111",
		01234 => "11111111",
		01235 => "11111111",
		01236 => "11111111",
		01237 => "11111111",
		01238 => "11111111",
		01239 => "11111111",
		01240 => "11111111",
		01241 => "11111111",
		01242 => "11111111",
		01243 => "11111111",
		01244 => "11111111",
		01245 => "11111111",
		01246 => "11111111",
		01247 => "11111111",
		01248 => "11111111",
		01249 => "11111111",
		01250 => "11111111",
		01251 => "11111111",
		01252 => "11111111",
		01253 => "11111111",
		01254 => "11111111",
		01255 => "11111111",
		01256 => "11111111",
		01257 => "11111111",
		01258 => "11111111",
		01259 => "11111111",
		01260 => "11111111",
		01261 => "11111111",
		01262 => "11111111",
		01263 => "11111111",
		01264 => "11111111",
		01265 => "11111111",
		01266 => "11111111",
		01267 => "11111111",
		01268 => "11111111",
		01269 => "11111111",
		01270 => "11111111",
		01271 => "11111111",
		01272 => "11111111",
		01273 => "11111111",
		01274 => "11111111",
		01275 => "11111111",
		01276 => "11111111",
		01277 => "11111111",
		01278 => "11111111",
		01279 => "11111111",
		01280 => "11111111",
		01281 => "11111111",
		01282 => "11111111",
		01283 => "11111111",
		01284 => "11111111",
		01285 => "11111111",
		01286 => "11111111",
		01287 => "11111111",
		01288 => "11111111",
		01289 => "11111111",
		01290 => "11111111",
		01291 => "11111111",
		01292 => "11111111",
		01293 => "11111111",
		01294 => "11111111",
		01295 => "11111111",
		01296 => "11111111",
		01297 => "11111111",
		01298 => "11111111",
		01299 => "11111111",
		01300 => "11111111",
		01301 => "11111111",
		01302 => "11111111",
		01303 => "11111111",
		01304 => "11111111",
		01305 => "11111111",
		01306 => "11111111",
		01307 => "11111111",
		01308 => "11111111",
		01309 => "11111111",
		01310 => "11111111",
		01311 => "11111111",
		01312 => "11111111",
		01313 => "11111111",
		01314 => "11111111",
		01315 => "11111111",
		01316 => "11111111",
		01317 => "11111111",
		01318 => "11111111",
		01319 => "11111111",
		01320 => "11111111",
		01321 => "11111111",
		01322 => "11111111",
		01323 => "11111111",
		01324 => "11111111",
		01325 => "11111111",
		01326 => "11111111",
		01327 => "11111111",
		01328 => "11111111",
		01329 => "11111111",
		01330 => "11111111",
		01331 => "11111111",
		01332 => "11111111",
		01333 => "11111111",
		01334 => "11111111",
		01335 => "11111111",
		01336 => "11111111",
		01337 => "11111111",
		01338 => "11111111",
		01339 => "11111111",
		01340 => "11111111",
		01341 => "11111111",
		01342 => "11111111",
		01343 => "11111111",
		01344 => "11111111",
		01345 => "11111111",
		01346 => "11111111",
		01347 => "11111111",
		01348 => "11111111",
		01349 => "11111111",
		01350 => "11111111",
		01351 => "11111111",
		01352 => "11111111",
		01353 => "11111111",
		01354 => "11111111",
		01355 => "11111111",
		01356 => "11111111",
		01357 => "11111111",
		01358 => "11111111",
		01359 => "11111111",
		01360 => "11111111",
		01361 => "11111111",
		01362 => "11111111",
		01363 => "11111111",
		01364 => "11111111",
		01365 => "11111111",
		01366 => "11111111",
		01367 => "11111111",
		01368 => "11111111",
		01369 => "11111111",
		01370 => "11111111",
		01371 => "11111111",
		01372 => "11111111",
		01373 => "11111111",
		01374 => "11111111",
		01375 => "11111111",
		01376 => "11111111",
		01377 => "11111111",
		01378 => "11111111",
		01379 => "11111111",
		01380 => "11111111",
		01381 => "11111111",
		01382 => "11111111",
		01383 => "11111111",
		01384 => "11111111",
		01385 => "11111111",
		01386 => "11111111",
		01387 => "11111111",
		01388 => "11111111",
		01389 => "11111111",
		01390 => "11111111",
		01391 => "11111111",
		01392 => "11111111",
		01393 => "11111111",
		01394 => "11111111",
		01395 => "11111111",
		01396 => "11111111",
		01397 => "11111111",
		01398 => "11111111",
		01399 => "11111111",
		01400 => "11111111",
		01401 => "11111111",
		01402 => "11111111",
		01403 => "11111111",
		01404 => "11111111",
		01405 => "11111111",
		01406 => "11111111",
		01407 => "11111111",
		01408 => "11111111",
		01409 => "11111111",
		01410 => "11111111",
		01411 => "11111111",
		01412 => "11111111",
		01413 => "11111111",
		01414 => "11111111",
		01415 => "11111111",
		01416 => "11111111",
		01417 => "11111111",
		01418 => "11111111",
		01419 => "11111111",
		01420 => "11111111",
		01421 => "11111111",
		01422 => "11111111",
		01423 => "11111111",
		01424 => "11111111",
		01425 => "11111111",
		01426 => "11111111",
		01427 => "11111111",
		01428 => "11111111",
		01429 => "11111111",
		01430 => "11111111",
		01431 => "11111111",
		01432 => "11111111",
		01433 => "11111111",
		01434 => "11111111",
		01435 => "11111111",
		01436 => "11111111",
		01437 => "11111111",
		01438 => "11111111",
		01439 => "11111111",
		01440 => "11111111",
		01441 => "11111111",
		01442 => "11111111",
		01443 => "11111111",
		01444 => "11111111",
		01445 => "11111111",
		01446 => "11111111",
		01447 => "11111111",
		01448 => "11111111",
		01449 => "11111111",
		01450 => "11111111",
		01451 => "11111111",
		01452 => "11111111",
		01453 => "11111111",
		01454 => "11111111",
		01455 => "11111111",
		01456 => "11111111",
		01457 => "11111111",
		01458 => "11111111",
		01459 => "11111111",
		01460 => "11111111",
		01461 => "11111111",
		01462 => "11111111",
		01463 => "11111111",
		01464 => "11111111",
		01465 => "11111111",
		01466 => "11111111",
		01467 => "11111111",
		01468 => "11111111",
		01469 => "11111111",
		01470 => "11111111",
		01471 => "11111111",
		01472 => "11111111",
		01473 => "11111111",
		01474 => "11111111",
		01475 => "11111111",
		01476 => "11111111",
		01477 => "11111111",
		01478 => "11111111",
		01479 => "11111111",
		01480 => "11111111",
		01481 => "11111111",
		01482 => "11111111",
		01483 => "11111111",
		01484 => "11111111",
		01485 => "11111111",
		01486 => "11111111",
		01487 => "11111111",
		01488 => "11111111",
		01489 => "11111111",
		01490 => "11111111",
		01491 => "11111111",
		01492 => "11111111",
		01493 => "11111111",
		01494 => "11111111",
		01495 => "11111111",
		01496 => "11111111",
		01497 => "11111111",
		01498 => "11111111",
		01499 => "11111111",
		01500 => "11111111",
		01501 => "11111111",
		01502 => "11111111",
		01503 => "11111111",
		01504 => "11111111",
		01505 => "11111111",
		01506 => "11111111",
		01507 => "11111111",
		01508 => "11111111",
		01509 => "11111111",
		01510 => "11111111",
		01511 => "11111111",
		01512 => "11111111",
		01513 => "11111111",
		01514 => "11111111",
		01515 => "11111111",
		01516 => "11111111",
		01517 => "11111111",
		01518 => "11111111",
		01519 => "11111111",
		01520 => "11111111",
		01521 => "11111111",
		01522 => "11111111",
		01523 => "11111111",
		01524 => "11111111",
		01525 => "11111111",
		01526 => "11111111",
		01527 => "11111111",
		01528 => "11111111",
		01529 => "11111111",
		01530 => "11111111",
		01531 => "11111111",
		01532 => "11111111",
		01533 => "11111111",
		01534 => "11111111",
		01535 => "11111111",
		01536 => "11111111",
		01537 => "11111111",
		01538 => "11111111",
		01539 => "11111111",
		01540 => "11111111",
		01541 => "11111111",
		01542 => "11111111",
		01543 => "11111111",
		01544 => "11111111",
		01545 => "11111111",
		01546 => "11111111",
		01547 => "11111111",
		01548 => "11111111",
		01549 => "11111111",
		01550 => "11111111",
		01551 => "11111111",
		01552 => "11111111",
		01553 => "11111111",
		01554 => "11111111",
		01555 => "11111111",
		01556 => "11111111",
		01557 => "11111111",
		01558 => "11111111",
		01559 => "11111111",
		01560 => "11111111",
		01561 => "11111111",
		01562 => "11111111",
		01563 => "11111111",
		01564 => "11111111",
		01565 => "11111111",
		01566 => "11111111",
		01567 => "11111111",
		01568 => "11111111",
		01569 => "11111111",
		01570 => "11111111",
		01571 => "11111111",
		01572 => "11111111",
		01573 => "11111111",
		01574 => "11111111",
		01575 => "11111111",
		01576 => "11111111",
		01577 => "11111111",
		01578 => "11111111",
		01579 => "11111111",
		01580 => "11111111",
		01581 => "11111111",
		01582 => "11111111",
		01583 => "11111111",
		01584 => "11111111",
		01585 => "11111111",
		01586 => "11111111",
		01587 => "11111111",
		01588 => "11111111",
		01589 => "11111111",
		01590 => "11111111",
		01591 => "11111111",
		01592 => "11111111",
		01593 => "11111111",
		01594 => "11111111",
		01595 => "11111111",
		01596 => "11111111",
		01597 => "11111111",
		01598 => "11111111",
		01599 => "11111111",
		01600 => "11111111",
		01601 => "11111111",
		01602 => "11111111",
		01603 => "11111111",
		01604 => "11111111",
		01605 => "11111111",
		01606 => "11111111",
		01607 => "11111111",
		01608 => "11111111",
		01609 => "11111111",
		01610 => "11111111",
		01611 => "11111111",
		01612 => "11111111",
		01613 => "11111111",
		01614 => "11111111",
		01615 => "11111111",
		01616 => "11111111",
		01617 => "11111111",
		01618 => "11111111",
		01619 => "11111111",
		01620 => "11111111",
		01621 => "11111111",
		01622 => "11111111",
		01623 => "11111111",
		01624 => "11111111",
		01625 => "11111111",
		01626 => "11111111",
		01627 => "11111111",
		01628 => "11111111",
		01629 => "11111111",
		01630 => "11111111",
		01631 => "11111111",
		01632 => "11111111",
		01633 => "11111111",
		01634 => "11111111",
		01635 => "11111111",
		01636 => "11111111",
		01637 => "11111111",
		01638 => "11111111",
		01639 => "11111111",
		01640 => "11111111",
		01641 => "11111111",
		01642 => "11111111",
		01643 => "11111111",
		01644 => "11111111",
		01645 => "11111111",
		01646 => "11111111",
		01647 => "11111111",
		01648 => "11111111",
		01649 => "11111111",
		01650 => "11111111",
		01651 => "11111111",
		01652 => "11111111",
		01653 => "11111111",
		01654 => "11111111",
		01655 => "11111111",
		01656 => "11111111",
		01657 => "11111111",
		01658 => "11111111",
		01659 => "11111111",
		01660 => "11111111",
		01661 => "11111111",
		01662 => "11111111",
		01663 => "11111111",
		01664 => "11111111",
		01665 => "11111111",
		01666 => "11111111",
		01667 => "11111111",
		01668 => "11111111",
		01669 => "11111111",
		01670 => "11111111",
		01671 => "11111111",
		01672 => "11111111",
		01673 => "11111111",
		01674 => "11111111",
		01675 => "11111111",
		01676 => "11111111",
		01677 => "11111111",
		01678 => "11111111",
		01679 => "11111111",
		01680 => "11111111",
		01681 => "11111111",
		01682 => "11111111",
		01683 => "11111111",
		01684 => "11111111",
		01685 => "11111111",
		01686 => "11111111",
		01687 => "11111111",
		01688 => "11111111",
		01689 => "11111111",
		01690 => "11111111",
		01691 => "11111111",
		01692 => "11111111",
		01693 => "11111111",
		01694 => "11111111",
		01695 => "11111111",
		01696 => "11111111",
		01697 => "11111111",
		01698 => "11111111",
		01699 => "11111111",
		01700 => "11111111",
		01701 => "11111111",
		01702 => "11111111",
		01703 => "11111111",
		01704 => "11111111",
		01705 => "11111111",
		01706 => "11111111",
		01707 => "11111111",
		01708 => "11111111",
		01709 => "11111111",
		01710 => "11111111",
		01711 => "11111111",
		01712 => "11111111",
		01713 => "11111111",
		01714 => "11111111",
		01715 => "11111111",
		01716 => "11111111",
		01717 => "11111111",
		01718 => "11111111",
		01719 => "11111111",
		01720 => "11111111",
		01721 => "11111111",
		01722 => "11111111",
		01723 => "11111111",
		01724 => "11111111",
		01725 => "11111111",
		01726 => "11111111",
		01727 => "11111111",
		01728 => "11111111",
		01729 => "11111111",
		01730 => "11111111",
		01731 => "11111111",
		01732 => "11111111",
		01733 => "11111111",
		01734 => "11111111",
		01735 => "11111111",
		01736 => "11111111",
		01737 => "11111111",
		01738 => "11111111",
		01739 => "11111111",
		01740 => "11111111",
		01741 => "11111111",
		01742 => "11111111",
		01743 => "11111111",
		01744 => "11111111",
		01745 => "11111111",
		01746 => "11111111",
		01747 => "11111111",
		01748 => "11111111",
		01749 => "11111111",
		01750 => "11111111",
		01751 => "11111111",
		01752 => "11111111",
		01753 => "11111111",
		01754 => "11111111",
		01755 => "11111111",
		01756 => "11111111",
		01757 => "11111111",
		01758 => "11111111",
		01759 => "11111111",
		01760 => "11111111",
		01761 => "11111111",
		01762 => "11111111",
		01763 => "11111111",
		01764 => "11111111",
		01765 => "11111111",
		01766 => "11111111",
		01767 => "11111111",
		01768 => "11111111",
		01769 => "11111111",
		01770 => "11111111",
		01771 => "11111111",
		01772 => "11111111",
		01773 => "11111111",
		01774 => "11111111",
		01775 => "11111111",
		01776 => "11111111",
		01777 => "11111111",
		01778 => "11111111",
		01779 => "11111111",
		01780 => "11111111",
		01781 => "11111111",
		01782 => "11111111",
		01783 => "11111111",
		01784 => "11111111",
		01785 => "11111111",
		01786 => "11111111",
		01787 => "11111111",
		01788 => "11111111",
		01789 => "11111111",
		01790 => "11111111",
		01791 => "11111111",
		01792 => "11111111",
		01793 => "11111111",
		01794 => "11111111",
		01795 => "11111111",
		01796 => "11111111",
		01797 => "11111111",
		01798 => "11111111",
		01799 => "11111111",
		01800 => "11111111",
		01801 => "11111111",
		01802 => "11111111",
		01803 => "11111111",
		01804 => "11111111",
		01805 => "11111111",
		01806 => "11111111",
		01807 => "11111111",
		01808 => "11111111",
		01809 => "11111111",
		01810 => "11111111",
		01811 => "11111111",
		01812 => "11111111",
		01813 => "11111111",
		01814 => "11111111",
		01815 => "11111111",
		01816 => "11111111",
		01817 => "11111111",
		01818 => "11111111",
		01819 => "11111111",
		01820 => "11111111",
		01821 => "11111111",
		01822 => "11111111",
		01823 => "11111111",
		01824 => "11111111",
		01825 => "11111111",
		01826 => "11111111",
		01827 => "11111111",
		01828 => "11111111",
		01829 => "11111111",
		01830 => "11111111",
		01831 => "11111111",
		01832 => "11111111",
		01833 => "11111111",
		01834 => "11111111",
		01835 => "11111111",
		01836 => "11111111",
		01837 => "11111111",
		01838 => "11111111",
		01839 => "11111111",
		01840 => "11111111",
		01841 => "11111111",
		01842 => "11111111",
		01843 => "11111111",
		01844 => "11111111",
		01845 => "11111111",
		01846 => "11111111",
		01847 => "11111111",
		01848 => "11111111",
		01849 => "11111111",
		01850 => "11111111",
		01851 => "11111111",
		01852 => "11111111",
		01853 => "11111111",
		01854 => "11111111",
		01855 => "11111111",
		01856 => "11111111",
		01857 => "11111111",
		01858 => "11111111",
		01859 => "11111111",
		01860 => "11111111",
		01861 => "11111111",
		01862 => "11111111",
		01863 => "11111111",
		01864 => "11111111",
		01865 => "11111111",
		01866 => "11111111",
		01867 => "11111111",
		01868 => "11111111",
		01869 => "11111111",
		01870 => "11111111",
		01871 => "11111111",
		01872 => "11111111",
		01873 => "11111111",
		01874 => "11111111",
		01875 => "11111111",
		01876 => "11111111",
		01877 => "11111111",
		01878 => "11111111",
		01879 => "11111111",
		01880 => "11111111",
		01881 => "11111111",
		01882 => "11111111",
		01883 => "11111111",
		01884 => "11111111",
		01885 => "11111111",
		01886 => "11111111",
		01887 => "11111111",
		01888 => "11111111",
		01889 => "11111111",
		01890 => "11111111",
		01891 => "11111111",
		01892 => "11111111",
		01893 => "11111111",
		01894 => "11111111",
		01895 => "11111111",
		01896 => "11111111",
		01897 => "11111111",
		01898 => "11111111",
		01899 => "11111111",
		01900 => "11111111",
		01901 => "11111111",
		01902 => "11111111",
		01903 => "11111111",
		01904 => "11111111",
		01905 => "11111111",
		01906 => "11111111",
		01907 => "11111111",
		01908 => "11111111",
		01909 => "11111111",
		01910 => "11111111",
		01911 => "11111111",
		01912 => "11111111",
		01913 => "11111111",
		01914 => "11111111",
		01915 => "11111111",
		01916 => "11111111",
		01917 => "11111111",
		01918 => "11111111",
		01919 => "11111111",
		01920 => "11111111",
		01921 => "11111111",
		01922 => "11111111",
		01923 => "11111111",
		01924 => "11111111",
		01925 => "11111111",
		01926 => "11111111",
		01927 => "11111111",
		01928 => "11111111",
		01929 => "11111111",
		01930 => "11111111",
		01931 => "11111111",
		01932 => "11111111",
		01933 => "11111111",
		01934 => "11111111",
		01935 => "11111111",
		01936 => "11111111",
		01937 => "11111111",
		01938 => "11111111",
		01939 => "11111111",
		01940 => "11111111",
		01941 => "11111111",
		01942 => "11111111",
		01943 => "11111111",
		01944 => "11111111",
		01945 => "11111111",
		01946 => "11111111",
		01947 => "11111111",
		01948 => "11111111",
		01949 => "11111111",
		01950 => "11111111",
		01951 => "11111111",
		01952 => "11111111",
		01953 => "11111111",
		01954 => "11111111",
		01955 => "11111111",
		01956 => "11111111",
		01957 => "11111111",
		01958 => "11111111",
		01959 => "11111111",
		01960 => "11111111",
		01961 => "11111111",
		01962 => "11111111",
		01963 => "11111111",
		01964 => "11111111",
		01965 => "11111111",
		01966 => "11111111",
		01967 => "11111111",
		01968 => "11111111",
		01969 => "11111111",
		01970 => "11111111",
		01971 => "11111111",
		01972 => "11111111",
		01973 => "11111111",
		01974 => "11111111",
		01975 => "11111111",
		01976 => "11111111",
		01977 => "11111111",
		01978 => "11111111",
		01979 => "11111111",
		01980 => "11111111",
		01981 => "11111111",
		01982 => "11111111",
		01983 => "11111111",
		01984 => "11111111",
		01985 => "11111111",
		01986 => "11111111",
		01987 => "11111111",
		01988 => "11111111",
		01989 => "11111111",
		01990 => "11111111",
		01991 => "11111111",
		01992 => "11111111",
		01993 => "11111111",
		01994 => "11111111",
		01995 => "11111111",
		01996 => "11111111",
		01997 => "11111111",
		01998 => "11111111",
		01999 => "11111111",
		02000 => "11111111",
		02001 => "11111111",
		02002 => "11111111",
		02003 => "11111111",
		02004 => "11111111",
		02005 => "11111111",
		02006 => "11111111",
		02007 => "11111111",
		02008 => "11111111",
		02009 => "11111111",
		02010 => "11111111",
		02011 => "11111111",
		02012 => "11111111",
		02013 => "11111111",
		02014 => "11111111",
		02015 => "11111111",
		02016 => "11111111",
		02017 => "11111111",
		02018 => "11111111",
		02019 => "11111111",
		02020 => "11111111",
		02021 => "11111111",
		02022 => "11111111",
		02023 => "11111111",
		02024 => "11111111",
		02025 => "11111111",
		02026 => "11111111",
		02027 => "11111111",
		02028 => "11111111",
		02029 => "11111111",
		02030 => "11111111",
		02031 => "11111111",
		02032 => "11111111",
		02033 => "11111111",
		02034 => "11111111",
		02035 => "11111111",
		02036 => "11111111",
		02037 => "11111111",
		02038 => "11111111",
		02039 => "11111111",
		02040 => "11111111",
		02041 => "11111111",
		02042 => "11111111",
		02043 => "11111111",
		02044 => "11111111",
		02045 => "11111111",
		02046 => "11111111",
		02047 => "11111111",
		02048 => "11111111",
		02049 => "11111111",
		02050 => "11111111",
		02051 => "11111111",
		02052 => "11111111",
		02053 => "11111111",
		02054 => "11111111",
		02055 => "11111111",
		02056 => "11111111",
		02057 => "11111111",
		02058 => "11111111",
		02059 => "11111111",
		02060 => "11111111",
		02061 => "11111111",
		02062 => "11111111",
		02063 => "11111111",
		02064 => "11111111",
		02065 => "11111111",
		02066 => "11111111",
		02067 => "11111111",
		02068 => "11111111",
		02069 => "11111111",
		02070 => "11111111",
		02071 => "11111111",
		02072 => "11111111",
		02073 => "11111111",
		02074 => "11111111",
		02075 => "11111111",
		02076 => "11111111",
		02077 => "11111111",
		02078 => "11111111",
		02079 => "11111111",
		02080 => "11111111",
		02081 => "11111111",
		02082 => "11111111",
		02083 => "11111111",
		02084 => "11111111",
		02085 => "11111111",
		02086 => "11111111",
		02087 => "11111111",
		02088 => "11111111",
		02089 => "11111111",
		02090 => "11111111",
		02091 => "11111111",
		02092 => "11111111",
		02093 => "11111111",
		02094 => "11111111",
		02095 => "11111111",
		02096 => "11111111",
		02097 => "11111111",
		02098 => "11111111",
		02099 => "11111111",
		02100 => "11111111",
		02101 => "11111111",
		02102 => "11111111",
		02103 => "11111111",
		02104 => "11111111",
		02105 => "11111111",
		02106 => "11111111",
		02107 => "11111111",
		02108 => "11111111",
		02109 => "11111111",
		02110 => "11111111",
		02111 => "11111111",
		02112 => "11111111",
		02113 => "11111111",
		02114 => "11111111",
		02115 => "11111111",
		02116 => "11111111",
		02117 => "11111111",
		02118 => "11111111",
		02119 => "11111111",
		02120 => "11111111",
		02121 => "11111111",
		02122 => "11111111",
		02123 => "11111111",
		02124 => "11111111",
		02125 => "11111111",
		02126 => "11111111",
		02127 => "11111111",
		02128 => "11111111",
		02129 => "11111111",
		02130 => "11111111",
		02131 => "11111111",
		02132 => "11111111",
		02133 => "11111111",
		02134 => "11111111",
		02135 => "11111111",
		02136 => "11111111",
		02137 => "11111111",
		02138 => "11111111",
		02139 => "11111111",
		02140 => "11111111",
		02141 => "11111111",
		02142 => "11111111",
		02143 => "11111111",
		02144 => "11111111",
		02145 => "11111111",
		02146 => "11111111",
		02147 => "11111111",
		02148 => "11111111",
		02149 => "11111111",
		02150 => "11111111",
		02151 => "11111111",
		02152 => "11111111",
		02153 => "11111111",
		02154 => "11111111",
		02155 => "11111111",
		02156 => "11111111",
		02157 => "11111111",
		02158 => "11111111",
		02159 => "11111111",
		02160 => "11111111",
		02161 => "11111111",
		02162 => "11111111",
		02163 => "11111111",
		02164 => "11111111",
		02165 => "11111111",
		02166 => "11111111",
		02167 => "11111111",
		02168 => "11111111",
		02169 => "11111111",
		02170 => "11111111",
		02171 => "11111111",
		02172 => "11111111",
		02173 => "11111111",
		02174 => "11111111",
		02175 => "11111111",
		02176 => "11111111",
		02177 => "11111111",
		02178 => "11111111",
		02179 => "11111111",
		02180 => "11111111",
		02181 => "11111111",
		02182 => "11111111",
		02183 => "11111111",
		02184 => "11111111",
		02185 => "11111111",
		02186 => "11111111",
		02187 => "11111111",
		02188 => "11111111",
		02189 => "11111111",
		02190 => "11111111",
		02191 => "11111111",
		02192 => "11111111",
		02193 => "11111111",
		02194 => "11111111",
		02195 => "11111111",
		02196 => "11111111",
		02197 => "11111111",
		02198 => "11111111",
		02199 => "11111111",
		02200 => "11111111",
		02201 => "11111111",
		02202 => "11111111",
		02203 => "11111111",
		02204 => "11111111",
		02205 => "11111111",
		02206 => "11111111",
		02207 => "11111111",
		02208 => "11111111",
		02209 => "11111111",
		02210 => "11111111",
		02211 => "11111111",
		02212 => "11111111",
		02213 => "11111111",
		02214 => "11111111",
		02215 => "11111111",
		02216 => "11111111",
		02217 => "11111111",
		02218 => "11111111",
		02219 => "11111111",
		02220 => "11111111",
		02221 => "11111111",
		02222 => "11111111",
		02223 => "11111111",
		02224 => "11111111",
		02225 => "11111111",
		02226 => "11111111",
		02227 => "11111111",
		02228 => "11111111",
		02229 => "11111111",
		02230 => "11111111",
		02231 => "11111111",
		02232 => "11111111",
		02233 => "11111111",
		02234 => "11111111",
		02235 => "11111111",
		02236 => "11111111",
		02237 => "11111111",
		02238 => "11111111",
		02239 => "11111111",
		02240 => "11111111",
		02241 => "11111111",
		02242 => "11111111",
		02243 => "11111111",
		02244 => "11111111",
		02245 => "11111111",
		02246 => "11111111",
		02247 => "11111111",
		02248 => "11111111",
		02249 => "11111111",
		02250 => "11111111",
		02251 => "11111111",
		02252 => "11111111",
		02253 => "11111111",
		02254 => "11111111",
		02255 => "11111111",
		02256 => "11111111",
		02257 => "11111111",
		02258 => "11111111",
		02259 => "11111111",
		02260 => "11111111",
		02261 => "11111111",
		02262 => "11111111",
		02263 => "11111111",
		02264 => "11111111",
		02265 => "11111111",
		02266 => "11111111",
		02267 => "11111111",
		02268 => "11111111",
		02269 => "11111111",
		02270 => "11111111",
		02271 => "11111111",
		02272 => "11111111",
		02273 => "11111111",
		02274 => "11111111",
		02275 => "11111111",
		02276 => "11111111",
		02277 => "11111111",
		02278 => "11111111",
		02279 => "11111111",
		02280 => "11111111",
		02281 => "11111111",
		02282 => "11111111",
		02283 => "11111111",
		02284 => "11111111",
		02285 => "11111111",
		02286 => "11111111",
		02287 => "11111111",
		02288 => "11111111",
		02289 => "11111111",
		02290 => "11111111",
		02291 => "11111111",
		02292 => "11111111",
		02293 => "11111111",
		02294 => "11111111",
		02295 => "11111111",
		02296 => "11111111",
		02297 => "11111111",
		02298 => "11111111",
		02299 => "11111111",
		02300 => "11111111",
		02301 => "11111111",
		02302 => "11111111",
		02303 => "11111111",
		02304 => "11111111",
		02305 => "11111111",
		02306 => "11111111",
		02307 => "11111111",
		02308 => "11111111",
		02309 => "11111111",
		02310 => "11111111",
		02311 => "11111111",
		02312 => "11111111",
		02313 => "11111111",
		02314 => "11111111",
		02315 => "11111111",
		02316 => "11111111",
		02317 => "11111111",
		02318 => "11111111",
		02319 => "11111111",
		02320 => "11111111",
		02321 => "11111111",
		02322 => "11111111",
		02323 => "11111111",
		02324 => "11111111",
		02325 => "11111111",
		02326 => "11111111",
		02327 => "11111111",
		02328 => "11111111",
		02329 => "11111111",
		02330 => "11111111",
		02331 => "11111111",
		02332 => "11111111",
		02333 => "11111111",
		02334 => "11111111",
		02335 => "11111111",
		02336 => "11111111",
		02337 => "11111111",
		02338 => "11111111",
		02339 => "11111111",
		02340 => "11111111",
		02341 => "11111111",
		02342 => "11111111",
		02343 => "11111111",
		02344 => "11111111",
		02345 => "11111111",
		02346 => "11111111",
		02347 => "11111111",
		02348 => "11111111",
		02349 => "11111111",
		02350 => "11111111",
		02351 => "11111111",
		02352 => "11111111",
		02353 => "11111111",
		02354 => "11111111",
		02355 => "11111111",
		02356 => "11111111",
		02357 => "11111111",
		02358 => "11111111",
		02359 => "11111111",
		02360 => "11111111",
		02361 => "11111111",
		02362 => "11111111",
		02363 => "11111111",
		02364 => "11111111",
		02365 => "11111111",
		02366 => "11111111",
		02367 => "11111111",
		02368 => "11111111",
		02369 => "11111111",
		02370 => "11111111",
		02371 => "11111111",
		02372 => "11111111",
		02373 => "11111111",
		02374 => "11111111",
		02375 => "11111111",
		02376 => "11111111",
		02377 => "11111111",
		02378 => "11111111",
		02379 => "11111111",
		02380 => "11111111",
		02381 => "11111111",
		02382 => "11111111",
		02383 => "11111111",
		02384 => "11111111",
		02385 => "11111111",
		02386 => "11111111",
		02387 => "11111111",
		02388 => "11111111",
		02389 => "11111111",
		02390 => "11111111",
		02391 => "11111111",
		02392 => "11111111",
		02393 => "11111111",
		02394 => "11111111",
		02395 => "11111111",
		02396 => "11111111",
		02397 => "11111111",
		02398 => "11111111",
		02399 => "11111111",
		02400 => "11111111",
		02401 => "11111111",
		02402 => "11111111",
		02403 => "11111111",
		02404 => "11111111",
		02405 => "11111111",
		02406 => "11111111",
		02407 => "11111111",
		02408 => "11111111",
		02409 => "11111111",
		02410 => "11111111",
		02411 => "11111111",
		02412 => "11111111",
		02413 => "11111111",
		02414 => "11111111",
		02415 => "11111111",
		02416 => "11111111",
		02417 => "11111111",
		02418 => "11111111",
		02419 => "11111111",
		02420 => "11111111",
		02421 => "11111111",
		02422 => "11111111",
		02423 => "11111111",
		02424 => "11111111",
		02425 => "11111111",
		02426 => "11111111",
		02427 => "11111111",
		02428 => "11111111",
		02429 => "11111111",
		02430 => "11111111",
		02431 => "11111111",
		02432 => "11111111",
		02433 => "11111111",
		02434 => "11111111",
		02435 => "11111111",
		02436 => "11111111",
		02437 => "11111111",
		02438 => "11111111",
		02439 => "11111111",
		02440 => "11111111",
		02441 => "11111111",
		02442 => "11111111",
		02443 => "11111111",
		02444 => "11111111",
		02445 => "11111111",
		02446 => "11111111",
		02447 => "11111111",
		02448 => "11111111",
		02449 => "11111111",
		02450 => "11111111",
		02451 => "11111111",
		02452 => "11111111",
		02453 => "11111111",
		02454 => "11111111",
		02455 => "11111111",
		02456 => "11111111",
		02457 => "11111111",
		02458 => "11111111",
		02459 => "11111111",
		02460 => "11111111",
		02461 => "11111111",
		02462 => "11111111",
		02463 => "11111111",
		02464 => "11111111",
		02465 => "11111111",
		02466 => "11111111",
		02467 => "11111111",
		02468 => "11111111",
		02469 => "11111111",
		02470 => "11111111",
		02471 => "11111111",
		02472 => "11111111",
		02473 => "11111111",
		02474 => "11111111",
		02475 => "11111111",
		02476 => "11111111",
		02477 => "11111111",
		02478 => "11111111",
		02479 => "11111111",
		02480 => "11111111",
		02481 => "11111111",
		02482 => "11111111",
		02483 => "11111111",
		02484 => "11111111",
		02485 => "11111111",
		02486 => "11111111",
		02487 => "11111111",
		02488 => "11111111",
		02489 => "11111111",
		02490 => "11111111",
		02491 => "11111111",
		02492 => "11111111",
		02493 => "11111111",
		02494 => "11111111",
		02495 => "11111111",
		02496 => "11111111",
		02497 => "11111111",
		02498 => "11111111",
		02499 => "11111111",
		02500 => "11111111",
		02501 => "11111111",
		02502 => "11111111",
		02503 => "11111111",
		02504 => "11111111",
		02505 => "11111111",
		02506 => "11111111",
		02507 => "11111111",
		02508 => "11111111",
		02509 => "11111111",
		02510 => "11111111",
		02511 => "11111111",
		02512 => "11111111",
		02513 => "11111111",
		02514 => "11111111",
		02515 => "11111111",
		02516 => "11111111",
		02517 => "11111111",
		02518 => "11111111",
		02519 => "11111111",
		02520 => "11111111",
		02521 => "11111111",
		02522 => "11111111",
		02523 => "11111111",
		02524 => "11111111",
		02525 => "11111111",
		02526 => "11111111",
		02527 => "11111111",
		02528 => "11111111",
		02529 => "11111111",
		02530 => "11111111",
		02531 => "11111111",
		02532 => "11111111",
		02533 => "11111111",
		02534 => "11111111",
		02535 => "11111111",
		02536 => "11111111",
		02537 => "11111111",
		02538 => "11111111",
		02539 => "11111111",
		02540 => "11111111",
		02541 => "11111111",
		02542 => "11111111",
		02543 => "11111111",
		02544 => "11111111",
		02545 => "11111111",
		02546 => "11111111",
		02547 => "11111111",
		02548 => "11111111",
		02549 => "11111111",
		02550 => "11111111",
		02551 => "11111111",
		02552 => "11111111",
		02553 => "11111111",
		02554 => "11111111",
		02555 => "11111111",
		02556 => "11111111",
		02557 => "11111111",
		02558 => "11111111",
		02559 => "11111111",
		02560 => "11111111",
		02561 => "11111111",
		02562 => "11111111",
		02563 => "11111111",
		02564 => "11111111",
		02565 => "11111111",
		02566 => "11111111",
		02567 => "11111111",
		02568 => "11111111",
		02569 => "11111111",
		02570 => "11111111",
		02571 => "11111111",
		02572 => "11111111",
		02573 => "11111111",
		02574 => "11111111",
		02575 => "11111111",
		02576 => "11111111",
		02577 => "11111111",
		02578 => "11111111",
		02579 => "11111111",
		02580 => "11111111",
		02581 => "11111111",
		02582 => "11111111",
		02583 => "11111111",
		02584 => "11111111",
		02585 => "11111111",
		02586 => "11111111",
		02587 => "11111111",
		02588 => "11111111",
		02589 => "11111111",
		02590 => "11111111",
		02591 => "11111111",
		02592 => "11111111",
		02593 => "11111111",
		02594 => "11111111",
		02595 => "11111111",
		02596 => "11111111",
		02597 => "11111111",
		02598 => "11111111",
		02599 => "11111111",
		02600 => "11111111",
		02601 => "11111111",
		02602 => "11111111",
		02603 => "11111111",
		02604 => "11111111",
		02605 => "11111111",
		02606 => "11111111",
		02607 => "11111111",
		02608 => "11111111",
		02609 => "11111111",
		02610 => "11111111",
		02611 => "11111111",
		02612 => "11111111",
		02613 => "11111111",
		02614 => "11111111",
		02615 => "11111111",
		02616 => "11111111",
		02617 => "11111111",
		02618 => "11111111",
		02619 => "11111111",
		02620 => "11111111",
		02621 => "11111111",
		02622 => "11111111",
		02623 => "11111111",
		02624 => "11111111",
		02625 => "11111111",
		02626 => "11111111",
		02627 => "11111111",
		02628 => "11111111",
		02629 => "11111111",
		02630 => "11111111",
		02631 => "11111111",
		02632 => "11111111",
		02633 => "11111111",
		02634 => "11111111",
		02635 => "11111111",
		02636 => "11111111",
		02637 => "11111111",
		02638 => "11111111",
		02639 => "11111111",
		02640 => "11111111",
		02641 => "11111111",
		02642 => "11111111",
		02643 => "11111111",
		02644 => "11111111",
		02645 => "11111111",
		02646 => "11111111",
		02647 => "11111111",
		02648 => "11111111",
		02649 => "11111111",
		02650 => "11111111",
		02651 => "11111111",
		02652 => "11111111",
		02653 => "11111111",
		02654 => "11111111",
		02655 => "11111111",
		02656 => "11111111",
		02657 => "11111111",
		02658 => "11111111",
		02659 => "11111111",
		02660 => "11111111",
		02661 => "11111111",
		02662 => "11111111",
		02663 => "11111111",
		02664 => "11111111",
		02665 => "11111111",
		02666 => "11111111",
		02667 => "11111111",
		02668 => "11111111",
		02669 => "11111111",
		02670 => "11111111",
		02671 => "11111111",
		02672 => "11111111",
		02673 => "11111111",
		02674 => "11111111",
		02675 => "11111111",
		02676 => "11111111",
		02677 => "11111111",
		02678 => "11111111",
		02679 => "11111111",
		02680 => "11111111",
		02681 => "11111111",
		02682 => "11111111",
		02683 => "11111111",
		02684 => "11111111",
		02685 => "11111111",
		02686 => "11111111",
		02687 => "11111111",
		02688 => "11111111",
		02689 => "11111111",
		02690 => "11111111",
		02691 => "11111111",
		02692 => "11111111",
		02693 => "11111111",
		02694 => "11111111",
		02695 => "11111111",
		02696 => "11111111",
		02697 => "11111111",
		02698 => "11111111",
		02699 => "11111111",
		02700 => "11111111",
		02701 => "11111111",
		02702 => "11111111",
		02703 => "11111111",
		02704 => "11111111",
		02705 => "11111111",
		02706 => "11111111",
		02707 => "11111111",
		02708 => "11111111",
		02709 => "11111111",
		02710 => "11111111",
		02711 => "11111111",
		02712 => "11111111",
		02713 => "11111111",
		02714 => "11111111",
		02715 => "11111111",
		02716 => "11111111",
		02717 => "11111111",
		02718 => "11111111",
		02719 => "11111111",
		02720 => "11111111",
		02721 => "11111111",
		02722 => "11111111",
		02723 => "11111111",
		02724 => "11111111",
		02725 => "11111111",
		02726 => "11111111",
		02727 => "11111111",
		02728 => "11111111",
		02729 => "11111111",
		02730 => "11111111",
		02731 => "11111111",
		02732 => "11111111",
		02733 => "11111111",
		02734 => "11111111",
		02735 => "11111111",
		02736 => "11111111",
		02737 => "11111111",
		02738 => "11111111",
		02739 => "11111111",
		02740 => "11111111",
		02741 => "11111111",
		02742 => "11111111",
		02743 => "11111111",
		02744 => "11111111",
		02745 => "11111111",
		02746 => "11111111",
		02747 => "11111111",
		02748 => "11111111",
		02749 => "11111111",
		02750 => "11111111",
		02751 => "11111111",
		02752 => "11111111",
		02753 => "11111111",
		02754 => "11111111",
		02755 => "11111111",
		02756 => "11111111",
		02757 => "11111111",
		02758 => "11111111",
		02759 => "11111111",
		02760 => "11111111",
		02761 => "11111111",
		02762 => "11111111",
		02763 => "11111111",
		02764 => "11111111",
		02765 => "11111111",
		02766 => "11111111",
		02767 => "11111111",
		02768 => "11111111",
		02769 => "11111111",
		02770 => "11111111",
		02771 => "11111111",
		02772 => "11111111",
		02773 => "11111111",
		02774 => "11111111",
		02775 => "11111111",
		02776 => "11111111",
		02777 => "11111111",
		02778 => "11111111",
		02779 => "11111111",
		02780 => "11111111",
		02781 => "11111111",
		02782 => "11111111",
		02783 => "11111111",
		02784 => "11111111",
		02785 => "11111111",
		02786 => "11111111",
		02787 => "11111111",
		02788 => "11111111",
		02789 => "11111111",
		02790 => "11111111",
		02791 => "11111111",
		02792 => "11111111",
		02793 => "11111111",
		02794 => "11111111",
		02795 => "11111111",
		02796 => "11111111",
		02797 => "11111111",
		02798 => "11111111",
		02799 => "11111111",
		02800 => "11111111",
		02801 => "11111111",
		02802 => "11111111",
		02803 => "11111111",
		02804 => "11111111",
		02805 => "11111111",
		02806 => "11111111",
		02807 => "11111111",
		02808 => "11111111",
		02809 => "11111111",
		02810 => "11111111",
		02811 => "11111111",
		02812 => "11111111",
		02813 => "11111111",
		02814 => "11111111",
		02815 => "11111111",
		02816 => "11111111",
		02817 => "11111111",
		02818 => "11111111",
		02819 => "11111111",
		02820 => "11111111",
		02821 => "11111111",
		02822 => "11111111",
		02823 => "11111111",
		02824 => "11111111",
		02825 => "11111111",
		02826 => "11111111",
		02827 => "11111111",
		02828 => "11111111",
		02829 => "11111111",
		02830 => "11111111",
		02831 => "11111111",
		02832 => "11111111",
		02833 => "11111111",
		02834 => "11111111",
		02835 => "11111111",
		02836 => "11111111",
		02837 => "11111111",
		02838 => "11111111",
		02839 => "11111111",
		02840 => "11111111",
		02841 => "11111111",
		02842 => "11111111",
		02843 => "11111111",
		02844 => "11111111",
		02845 => "11111111",
		02846 => "11111111",
		02847 => "11111111",
		02848 => "11111111",
		02849 => "11111111",
		02850 => "11111111",
		02851 => "11111111",
		02852 => "11111111",
		02853 => "11111111",
		02854 => "11111111",
		02855 => "11111111",
		02856 => "11111111",
		02857 => "11111111",
		02858 => "11111111",
		02859 => "11111111",
		02860 => "11111111",
		02861 => "11111111",
		02862 => "11111111",
		02863 => "11111111",
		02864 => "11111111",
		02865 => "11111111",
		02866 => "11111111",
		02867 => "11111111",
		02868 => "11111111",
		02869 => "11111111",
		02870 => "11111111",
		02871 => "11111111",
		02872 => "11111111",
		02873 => "11111111",
		02874 => "11111111",
		02875 => "11111111",
		02876 => "11111111",
		02877 => "11111111",
		02878 => "11111111",
		02879 => "11111111",
		02880 => "11111111",
		02881 => "11111111",
		02882 => "11111111",
		02883 => "11111111",
		02884 => "11111111",
		02885 => "11111111",
		02886 => "11111111",
		02887 => "11111111",
		02888 => "11111111",
		02889 => "11111111",
		02890 => "11111111",
		02891 => "11111111",
		02892 => "11111111",
		02893 => "11111111",
		02894 => "11111111",
		02895 => "11111111",
		02896 => "11111111",
		02897 => "11111111",
		02898 => "11111111",
		02899 => "11111111",
		02900 => "11111111",
		02901 => "11111111",
		02902 => "11111111",
		02903 => "11111111",
		02904 => "11111111",
		02905 => "11111111",
		02906 => "11111111",
		02907 => "11111111",
		02908 => "11111111",
		02909 => "11111111",
		02910 => "11111111",
		02911 => "11111111",
		02912 => "11111111",
		02913 => "11111111",
		02914 => "11111111",
		02915 => "11111111",
		02916 => "11111111",
		02917 => "11111111",
		02918 => "11111111",
		02919 => "11111111",
		02920 => "11111111",
		02921 => "11111111",
		02922 => "11111111",
		02923 => "11111111",
		02924 => "11111111",
		02925 => "11111111",
		02926 => "11111111",
		02927 => "11111111",
		02928 => "11111111",
		02929 => "11111111",
		02930 => "11111111",
		02931 => "11111111",
		02932 => "11111111",
		02933 => "11111111",
		02934 => "11111111",
		02935 => "11111111",
		02936 => "11111111",
		02937 => "11111111",
		02938 => "11111111",
		02939 => "11111111",
		02940 => "11111111",
		02941 => "11111111",
		02942 => "11111111",
		02943 => "11111111",
		02944 => "11111111",
		02945 => "11111111",
		02946 => "11111111",
		02947 => "11111111",
		02948 => "11111111",
		02949 => "11111111",
		02950 => "11111111",
		02951 => "11111111",
		02952 => "11111111",
		02953 => "11111111",
		02954 => "11111111",
		02955 => "11111111",
		02956 => "11111111",
		02957 => "11111111",
		02958 => "11111111",
		02959 => "11111111",
		02960 => "11111111",
		02961 => "11111111",
		02962 => "11111111",
		02963 => "11111111",
		02964 => "11111111",
		02965 => "11111111",
		02966 => "11111111",
		02967 => "11111111",
		02968 => "11111111",
		02969 => "11111111",
		02970 => "11111111",
		02971 => "11111111",
		02972 => "11111111",
		02973 => "11111111",
		02974 => "11111111",
		02975 => "11111111",
		02976 => "11111111",
		02977 => "11111111",
		02978 => "11111111",
		02979 => "11111111",
		02980 => "11111111",
		02981 => "11111111",
		02982 => "11111111",
		02983 => "11111111",
		02984 => "11111111",
		02985 => "11111111",
		02986 => "11111111",
		02987 => "11111111",
		02988 => "11111111",
		02989 => "11111111",
		02990 => "11111111",
		02991 => "11111111",
		02992 => "11111111",
		02993 => "11111111",
		02994 => "11111111",
		02995 => "11111111",
		02996 => "11111111",
		02997 => "11111111",
		02998 => "11111111",
		02999 => "11111111",
		03000 => "11111111",
		03001 => "11111111",
		03002 => "11111111",
		03003 => "11111111",
		03004 => "11111111",
		03005 => "11111111",
		03006 => "11111111",
		03007 => "11111111",
		03008 => "11111111",
		03009 => "11111111",
		03010 => "11111111",
		03011 => "11111111",
		03012 => "11111111",
		03013 => "11111111",
		03014 => "11111111",
		03015 => "11111111",
		03016 => "11111111",
		03017 => "11111111",
		03018 => "11111111",
		03019 => "11111111",
		03020 => "11111111",
		03021 => "11111111",
		03022 => "11111111",
		03023 => "11111111",
		03024 => "11111111",
		03025 => "11111111",
		03026 => "11111111",
		03027 => "11111111",
		03028 => "11111111",
		03029 => "11111111",
		03030 => "11111111",
		03031 => "11111111",
		03032 => "11111111",
		03033 => "11111111",
		03034 => "11111111",
		03035 => "11111111",
		03036 => "11111111",
		03037 => "11111111",
		03038 => "11111111",
		03039 => "11111111",
		03040 => "11111111",
		03041 => "11111111",
		03042 => "11111111",
		03043 => "11111111",
		03044 => "11111111",
		03045 => "11111111",
		03046 => "11111111",
		03047 => "11111111",
		03048 => "11111111",
		03049 => "11111111",
		03050 => "11111111",
		03051 => "11111111",
		03052 => "11111111",
		03053 => "11111111",
		03054 => "11111111",
		03055 => "11111111",
		03056 => "11111111",
		03057 => "11111111",
		03058 => "11111111",
		03059 => "11111111",
		03060 => "11111111",
		03061 => "11111111",
		03062 => "11111111",
		03063 => "11111111",
		03064 => "11111111",
		03065 => "11111111",
		03066 => "11111111",
		03067 => "11111111",
		03068 => "11111111",
		03069 => "11111111",
		03070 => "11111111",
		03071 => "11111111",
		03072 => "11111111",
		03073 => "11111111",
		03074 => "11111111",
		03075 => "11111111",
		03076 => "11111111",
		03077 => "11111111",
		03078 => "11111111",
		03079 => "11111111",
		03080 => "11111111",
		03081 => "11111111",
		03082 => "11111111",
		03083 => "11111111",
		03084 => "11111111",
		03085 => "11111111",
		03086 => "11111111",
		03087 => "11111111",
		03088 => "11111111",
		03089 => "11111111",
		03090 => "11111111",
		03091 => "11111111",
		03092 => "11111111",
		03093 => "11111111",
		03094 => "11111111",
		03095 => "11111111",
		03096 => "11111111",
		03097 => "11111111",
		03098 => "11111111",
		03099 => "11111111",
		03100 => "11111111",
		03101 => "11111111",
		03102 => "11111111",
		03103 => "11111111",
		03104 => "11111111",
		03105 => "11111111",
		03106 => "11111111",
		03107 => "11111111",
		03108 => "11111111",
		03109 => "11111111",
		03110 => "11111111",
		03111 => "11111111",
		03112 => "11111111",
		03113 => "11111111",
		03114 => "11111111",
		03115 => "11111111",
		03116 => "11111111",
		03117 => "11111111",
		03118 => "11111111",
		03119 => "11111111",
		03120 => "11111111",
		03121 => "11111111",
		03122 => "11111111",
		03123 => "11111111",
		03124 => "11111111",
		03125 => "11111111",
		03126 => "11111111",
		03127 => "11111111",
		03128 => "11111111",
		03129 => "11111111",
		03130 => "11111111",
		03131 => "11111111",
		03132 => "11111111",
		03133 => "11111111",
		03134 => "11111111",
		03135 => "11111111",
		03136 => "11111111",
		03137 => "11111111",
		03138 => "11111111",
		03139 => "11111111",
		03140 => "11111111",
		03141 => "11111111",
		03142 => "11111111",
		03143 => "11111111",
		03144 => "11111111",
		03145 => "11111111",
		03146 => "11111111",
		03147 => "11111111",
		03148 => "11111111",
		03149 => "11111111",
		03150 => "11111111",
		03151 => "11111111",
		03152 => "11111111",
		03153 => "11111111",
		03154 => "11111111",
		03155 => "11111111",
		03156 => "11111111",
		03157 => "11111111",
		03158 => "11111111",
		03159 => "11111111",
		03160 => "11111111",
		03161 => "11111111",
		03162 => "11111111",
		03163 => "11111111",
		03164 => "11111111",
		03165 => "11111111",
		03166 => "11111111",
		03167 => "11111111",
		03168 => "11111111",
		03169 => "11111111",
		03170 => "11111111",
		03171 => "11111111",
		03172 => "11111111",
		03173 => "11111111",
		03174 => "11111111",
		03175 => "11111111",
		03176 => "11111111",
		03177 => "11111111",
		03178 => "11111111",
		03179 => "11111111",
		03180 => "11111111",
		03181 => "11111111",
		03182 => "11111111",
		03183 => "11111111",
		03184 => "11111111",
		03185 => "11111111",
		03186 => "11111111",
		03187 => "11111111",
		03188 => "11111111",
		03189 => "11111111",
		03190 => "11111111",
		03191 => "11111111",
		03192 => "11111111",
		03193 => "11111111",
		03194 => "11111111",
		03195 => "11111111",
		03196 => "11111111",
		03197 => "11111111",
		03198 => "11111111",
		03199 => "11111111",
		03200 => "11111111",
		03201 => "11111111",
		03202 => "11111111",
		03203 => "11111111",
		03204 => "11111111",
		03205 => "11111111",
		03206 => "11111111",
		03207 => "11111111",
		03208 => "11111111",
		03209 => "11111111",
		03210 => "11111111",
		03211 => "11111111",
		03212 => "11111111",
		03213 => "11111111",
		03214 => "11111111",
		03215 => "11111111",
		03216 => "11111111",
		03217 => "11111111",
		03218 => "11111111",
		03219 => "11111111",
		03220 => "11111111",
		03221 => "11111111",
		03222 => "11111111",
		03223 => "11111111",
		03224 => "11111111",
		03225 => "11111111",
		03226 => "11111111",
		03227 => "11111111",
		03228 => "11111111",
		03229 => "11111111",
		03230 => "11111111",
		03231 => "11111111",
		03232 => "11111111",
		03233 => "11111111",
		03234 => "11111111",
		03235 => "11111111",
		03236 => "11111111",
		03237 => "11111111",
		03238 => "11111111",
		03239 => "11111111",
		03240 => "11111111",
		03241 => "11111111",
		03242 => "11111111",
		03243 => "11111111",
		03244 => "11111111",
		03245 => "11111111",
		03246 => "11111111",
		03247 => "11111111",
		03248 => "11111111",
		03249 => "11111111",
		03250 => "11111111",
		03251 => "11111111",
		03252 => "11111111",
		03253 => "11111111",
		03254 => "11111111",
		03255 => "11111111",
		03256 => "11111111",
		03257 => "11111111",
		03258 => "11111111",
		03259 => "11111111",
		03260 => "11111111",
		03261 => "11111111",
		03262 => "11111111",
		03263 => "11111111",
		03264 => "11111111",
		03265 => "11111111",
		03266 => "11111111",
		03267 => "11111111",
		03268 => "11111111",
		03269 => "11111111",
		03270 => "11111111",
		03271 => "11111111",
		03272 => "11111111",
		03273 => "11111111",
		03274 => "11111111",
		03275 => "11111111",
		03276 => "11111111",
		03277 => "11111111",
		03278 => "11111111",
		03279 => "11111111",
		03280 => "11111111",
		03281 => "11111111",
		03282 => "11111111",
		03283 => "11111111",
		03284 => "11111111",
		03285 => "11111111",
		03286 => "11111111",
		03287 => "11111111",
		03288 => "11111111",
		03289 => "11111111",
		03290 => "11111111",
		03291 => "11111111",
		03292 => "11111111",
		03293 => "11111111",
		03294 => "11111111",
		03295 => "11111111",
		03296 => "11111111",
		03297 => "11111111",
		03298 => "11111111",
		03299 => "11111111",
		03300 => "11111111",
		03301 => "11111111",
		03302 => "11111111",
		03303 => "11111111",
		03304 => "11111111",
		03305 => "11111111",
		03306 => "11111111",
		03307 => "11111111",
		03308 => "11111111",
		03309 => "11111111",
		03310 => "11111111",
		03311 => "11111111",
		03312 => "11111111",
		03313 => "11111111",
		03314 => "11111111",
		03315 => "11111111",
		03316 => "11111111",
		03317 => "11111111",
		03318 => "11111111",
		03319 => "11111111",
		03320 => "11111111",
		03321 => "11111111",
		03322 => "11111111",
		03323 => "11111111",
		03324 => "11111111",
		03325 => "11111111",
		03326 => "11111111",
		03327 => "11111111",
		03328 => "11111111",
		03329 => "11111111",
		03330 => "11111111",
		03331 => "11111111",
		03332 => "11111111",
		03333 => "11111111",
		03334 => "11111111",
		03335 => "11111111",
		03336 => "11111111",
		03337 => "11111111",
		03338 => "11111111",
		03339 => "11111111",
		03340 => "11111111",
		03341 => "11111111",
		03342 => "11111111",
		03343 => "11111111",
		03344 => "11111111",
		03345 => "11111111",
		03346 => "11111111",
		03347 => "11111111",
		03348 => "11111111",
		03349 => "11111111",
		03350 => "11111111",
		03351 => "11111111",
		03352 => "11111111",
		03353 => "11111111",
		03354 => "11111111",
		03355 => "11111111",
		03356 => "11111111",
		03357 => "11111111",
		03358 => "11111111",
		03359 => "11111111",
		03360 => "11111111",
		03361 => "11111111",
		03362 => "11111111",
		03363 => "11111111",
		03364 => "11111111",
		03365 => "11111111",
		03366 => "11111111",
		03367 => "11111111",
		03368 => "11111111",
		03369 => "11111111",
		03370 => "11111111",
		03371 => "11111111",
		03372 => "11111111",
		03373 => "11111111",
		03374 => "11111111",
		03375 => "11111111",
		03376 => "11111111",
		03377 => "11111111",
		03378 => "11111111",
		03379 => "11111111",
		03380 => "11111111",
		03381 => "11111111",
		03382 => "11111111",
		03383 => "11111111",
		03384 => "11111111",
		03385 => "11111111",
		03386 => "11111111",
		03387 => "11111111",
		03388 => "11111111",
		03389 => "11111111",
		03390 => "11111111",
		03391 => "11111111",
		03392 => "11111111",
		03393 => "11111111",
		03394 => "11111111",
		03395 => "11111111",
		03396 => "11111111",
		03397 => "11111111",
		03398 => "11111111",
		03399 => "11111111",
		03400 => "11111111",
		03401 => "11111111",
		03402 => "11111111",
		03403 => "11111111",
		03404 => "11111111",
		03405 => "11111111",
		03406 => "11111111",
		03407 => "11111111",
		03408 => "11111111",
		03409 => "11111111",
		03410 => "11111111",
		03411 => "11111111",
		03412 => "11111111",
		03413 => "11111111",
		03414 => "11111111",
		03415 => "11111111",
		03416 => "11111111",
		03417 => "11111111",
		03418 => "11111111",
		03419 => "11111111",
		03420 => "11111111",
		03421 => "11111111",
		03422 => "11111111",
		03423 => "11111111",
		03424 => "11111111",
		03425 => "11111111",
		03426 => "11111111",
		03427 => "11111111",
		03428 => "11111111",
		03429 => "11111111",
		03430 => "11111111",
		03431 => "11111111",
		03432 => "11111111",
		03433 => "11111111",
		03434 => "11111111",
		03435 => "11111111",
		03436 => "11111111",
		03437 => "11111111",
		03438 => "11111111",
		03439 => "11111111",
		03440 => "11111111",
		03441 => "11111111",
		03442 => "11111111",
		03443 => "11111111",
		03444 => "11111111",
		03445 => "11111111",
		03446 => "11111111",
		03447 => "11111111",
		03448 => "11111111",
		03449 => "11111111",
		03450 => "11111111",
		03451 => "11111111",
		03452 => "11111111",
		03453 => "11111111",
		03454 => "11111111",
		03455 => "11111111",
		03456 => "11111111",
		03457 => "11111111",
		03458 => "11111111",
		03459 => "11111111",
		03460 => "11111111",
		03461 => "11111111",
		03462 => "11111111",
		03463 => "11111111",
		03464 => "11111111",
		03465 => "11111111",
		03466 => "11111111",
		03467 => "11111111",
		03468 => "11111111",
		03469 => "11111111",
		03470 => "11111111",
		03471 => "11111111",
		03472 => "11111111",
		03473 => "11111111",
		03474 => "11111111",
		03475 => "11111111",
		03476 => "11111111",
		03477 => "11111111",
		03478 => "11111111",
		03479 => "11111111",
		03480 => "11111111",
		03481 => "11111111",
		03482 => "11111111",
		03483 => "11111111",
		03484 => "11111111",
		03485 => "11111111",
		03486 => "11111111",
		03487 => "11111111",
		03488 => "11111111",
		03489 => "11111111",
		03490 => "11111111",
		03491 => "11111111",
		03492 => "11111111",
		03493 => "11111111",
		03494 => "11111111",
		03495 => "11111111",
		03496 => "11111111",
		03497 => "11111111",
		03498 => "11111111",
		03499 => "11111111",
		03500 => "11111111",
		03501 => "11111111",
		03502 => "11111111",
		03503 => "11111111",
		03504 => "11111111",
		03505 => "11111111",
		03506 => "11111111",
		03507 => "11111111",
		03508 => "11111111",
		03509 => "11111111",
		03510 => "11111111",
		03511 => "11111111",
		03512 => "11111111",
		03513 => "11111111",
		03514 => "11111111",
		03515 => "11111111",
		03516 => "11111111",
		03517 => "11111111",
		03518 => "11111111",
		03519 => "11111111",
		03520 => "11111111",
		03521 => "11111111",
		03522 => "11111111",
		03523 => "11111111",
		03524 => "11111111",
		03525 => "11111111",
		03526 => "11111111",
		03527 => "11111111",
		03528 => "11111111",
		03529 => "11111111",
		03530 => "11111111",
		03531 => "11111111",
		03532 => "11111111",
		03533 => "11111111",
		03534 => "11111111",
		03535 => "11111111",
		03536 => "11111111",
		03537 => "11111111",
		03538 => "11111111",
		03539 => "11111111",
		03540 => "11111111",
		03541 => "11111111",
		03542 => "11111111",
		03543 => "11111111",
		03544 => "11111111",
		03545 => "11111111",
		03546 => "11111111",
		03547 => "11111111",
		03548 => "11111111",
		03549 => "11111111",
		03550 => "11111111",
		03551 => "11111111",
		03552 => "11111111",
		03553 => "11111111",
		03554 => "11111111",
		03555 => "11111111",
		03556 => "11111111",
		03557 => "11111111",
		03558 => "11111111",
		03559 => "11111111",
		03560 => "11111111",
		03561 => "11111111",
		03562 => "11111111",
		03563 => "11111111",
		03564 => "11111111",
		03565 => "11111111",
		03566 => "11111111",
		03567 => "11111111",
		03568 => "11111111",
		03569 => "11111111",
		03570 => "11111111",
		03571 => "11111111",
		03572 => "11111111",
		03573 => "11111111",
		03574 => "11111111",
		03575 => "11111111",
		03576 => "11111111",
		03577 => "11111111",
		03578 => "11111111",
		03579 => "11111111",
		03580 => "11111111",
		03581 => "11111111",
		03582 => "11111111",
		03583 => "11111111",
		03584 => "11111111",
		03585 => "11111111",
		03586 => "11111111",
		03587 => "11111111",
		03588 => "11111111",
		03589 => "11111111",
		03590 => "11111111",
		03591 => "11111111",
		03592 => "11111111",
		03593 => "11111111",
		03594 => "11111111",
		03595 => "11111111",
		03596 => "11111111",
		03597 => "11111111",
		03598 => "11111111",
		03599 => "11111111",
		03600 => "11111111",
		03601 => "11111111",
		03602 => "11111111",
		03603 => "11111111",
		03604 => "11111111",
		03605 => "11111111",
		03606 => "11111111",
		03607 => "11111111",
		03608 => "11111111",
		03609 => "11111111",
		03610 => "11111111",
		03611 => "11111111",
		03612 => "11111111",
		03613 => "11111111",
		03614 => "11111111",
		03615 => "11111111",
		03616 => "11111111",
		03617 => "11111111",
		03618 => "11111111",
		03619 => "11111111",
		03620 => "11111111",
		03621 => "11111111",
		03622 => "11111111",
		03623 => "11111111",
		03624 => "11111111",
		03625 => "11111111",
		03626 => "11111111",
		03627 => "11111111",
		03628 => "11111111",
		03629 => "11111111",
		03630 => "11111111",
		03631 => "11111111",
		03632 => "11111111",
		03633 => "11111111",
		03634 => "11111111",
		03635 => "11111111",
		03636 => "11111111",
		03637 => "11111111",
		03638 => "11111111",
		03639 => "11111111",
		03640 => "11111111",
		03641 => "11111111",
		03642 => "11111111",
		03643 => "11111111",
		03644 => "11111111",
		03645 => "11111111",
		03646 => "11111111",
		03647 => "11111111",
		03648 => "11111111",
		03649 => "11111111",
		03650 => "11111111",
		03651 => "11111111",
		03652 => "11111111",
		03653 => "11111111",
		03654 => "11111111",
		03655 => "11111111",
		03656 => "11111111",
		03657 => "11111111",
		03658 => "11111111",
		03659 => "11111111",
		03660 => "11111111",
		03661 => "11111111",
		03662 => "11111111",
		03663 => "11111111",
		03664 => "11111111",
		03665 => "11111111",
		03666 => "11111111",
		03667 => "11111111",
		03668 => "11111111",
		03669 => "11111111",
		03670 => "11111111",
		03671 => "11111111",
		03672 => "11111111",
		03673 => "11111111",
		03674 => "11111111",
		03675 => "11111111",
		03676 => "11111111",
		03677 => "11111111",
		03678 => "11111111",
		03679 => "11111111",
		03680 => "11111111",
		03681 => "11111111",
		03682 => "11111111",
		03683 => "11111111",
		03684 => "11111111",
		03685 => "11111111",
		03686 => "11111111",
		03687 => "11111111",
		03688 => "11111111",
		03689 => "11111111",
		03690 => "11111111",
		03691 => "11111111",
		03692 => "11111111",
		03693 => "11111111",
		03694 => "11111111",
		03695 => "11111111",
		03696 => "11111111",
		03697 => "11111111",
		03698 => "11111111",
		03699 => "11111111",
		03700 => "11111111",
		03701 => "11111111",
		03702 => "11111111",
		03703 => "11111111",
		03704 => "11111111",
		03705 => "11111111",
		03706 => "11111111",
		03707 => "11111111",
		03708 => "11111111",
		03709 => "11111111",
		03710 => "11111111",
		03711 => "11111111",
		03712 => "11111111",
		03713 => "11111111",
		03714 => "11111111",
		03715 => "11111111",
		03716 => "11111111",
		03717 => "11111111",
		03718 => "11111111",
		03719 => "11111111",
		03720 => "11111111",
		03721 => "11111111",
		03722 => "11111111",
		03723 => "11111111",
		03724 => "11111111",
		03725 => "11111111",
		03726 => "11111111",
		03727 => "11111111",
		03728 => "11111111",
		03729 => "11111111",
		03730 => "11111111",
		03731 => "11111111",
		03732 => "11111111",
		03733 => "11111111",
		03734 => "11111111",
		03735 => "11111111",
		03736 => "11111111",
		03737 => "11111111",
		03738 => "11111111",
		03739 => "11111111",
		03740 => "11111111",
		03741 => "11111111",
		03742 => "11111111",
		03743 => "11111111",
		03744 => "11111111",
		03745 => "11111111",
		03746 => "11111111",
		03747 => "11111111",
		03748 => "11111111",
		03749 => "11111111",
		03750 => "11111111",
		03751 => "11111111",
		03752 => "11111111",
		03753 => "11111111",
		03754 => "11111111",
		03755 => "11111111",
		03756 => "11111111",
		03757 => "11111111",
		03758 => "11111111",
		03759 => "11111111",
		03760 => "11111111",
		03761 => "11111111",
		03762 => "11111111",
		03763 => "11111111",
		03764 => "11111111",
		03765 => "11111111",
		03766 => "11111111",
		03767 => "11111111",
		03768 => "11111111",
		03769 => "11111111",
		03770 => "11111111",
		03771 => "11111111",
		03772 => "11111111",
		03773 => "11111111",
		03774 => "11111111",
		03775 => "11111111",
		03776 => "11111111",
		03777 => "11111111",
		03778 => "11111111",
		03779 => "11111111",
		03780 => "11111111",
		03781 => "11111111",
		03782 => "11111111",
		03783 => "11111111",
		03784 => "11111111",
		03785 => "11111111",
		03786 => "11111111",
		03787 => "11111111",
		03788 => "11111111",
		03789 => "11111111",
		03790 => "11111111",
		03791 => "11111111",
		03792 => "11111111",
		03793 => "11111111",
		03794 => "11111111",
		03795 => "11111111",
		03796 => "11111111",
		03797 => "11111111",
		03798 => "11111111",
		03799 => "11111111",
		03800 => "11111111",
		03801 => "11111111",
		03802 => "11111111",
		03803 => "11111111",
		03804 => "11111111",
		03805 => "11111111",
		03806 => "11111111",
		03807 => "11111111",
		03808 => "11111111",
		03809 => "11111111",
		03810 => "11111111",
		03811 => "11111111",
		03812 => "11111111",
		03813 => "11111111",
		03814 => "11111111",
		03815 => "11111111",
		03816 => "11111111",
		03817 => "11111111",
		03818 => "11111111",
		03819 => "11111111",
		03820 => "11111111",
		03821 => "11111111",
		03822 => "11111111",
		03823 => "11111111",
		03824 => "11111111",
		03825 => "11111111",
		03826 => "11111111",
		03827 => "11111111",
		03828 => "11111111",
		03829 => "11111111",
		03830 => "11111111",
		03831 => "11111111",
		03832 => "11111111",
		03833 => "11111111",
		03834 => "11111111",
		03835 => "11111111",
		03836 => "11111111",
		03837 => "11111111",
		03838 => "11111111",
		03839 => "11111111",
		03840 => "11111111",
		03841 => "11111111",
		03842 => "11111111",
		03843 => "11111111",
		03844 => "11111111",
		03845 => "11111111",
		03846 => "11111111",
		03847 => "11111111",
		03848 => "11111111",
		03849 => "11111111",
		03850 => "11111111",
		03851 => "11111111",
		03852 => "11111111",
		03853 => "11111111",
		03854 => "11111111",
		03855 => "11111111",
		03856 => "11111111",
		03857 => "11111111",
		03858 => "11111111",
		03859 => "11111111",
		03860 => "11111111",
		03861 => "11111111",
		03862 => "11111111",
		03863 => "11111111",
		03864 => "11111111",
		03865 => "11111111",
		03866 => "11111111",
		03867 => "11111111",
		03868 => "11111111",
		03869 => "11111111",
		03870 => "11111111",
		03871 => "11111111",
		03872 => "11111111",
		03873 => "11111111",
		03874 => "11111111",
		03875 => "11111111",
		03876 => "11111111",
		03877 => "11111111",
		03878 => "11111111",
		03879 => "11111111",
		03880 => "11111111",
		03881 => "11111111",
		03882 => "11111111",
		03883 => "11111111",
		03884 => "11111111",
		03885 => "11111111",
		03886 => "11111111",
		03887 => "11111111",
		03888 => "11111111",
		03889 => "11111111",
		03890 => "11111111",
		03891 => "11111111",
		03892 => "11111111",
		03893 => "11111111",
		03894 => "11111111",
		03895 => "11111111",
		03896 => "11111111",
		03897 => "11111111",
		03898 => "11111111",
		03899 => "11111111",
		03900 => "11111111",
		03901 => "11111111",
		03902 => "11111111",
		03903 => "11111111",
		03904 => "11111111",
		03905 => "11111111",
		03906 => "11111111",
		03907 => "11111111",
		03908 => "11111111",
		03909 => "11111111",
		03910 => "11111111",
		03911 => "11111111",
		03912 => "11111111",
		03913 => "11111111",
		03914 => "11111111",
		03915 => "11111111",
		03916 => "11111111",
		03917 => "11111111",
		03918 => "11111111",
		03919 => "11111111",
		03920 => "11111111",
		03921 => "11111111",
		03922 => "11111111",
		03923 => "11111111",
		03924 => "11111111",
		03925 => "11111111",
		03926 => "11111111",
		03927 => "11111111",
		03928 => "11111111",
		03929 => "11111111",
		03930 => "11111111",
		03931 => "11111111",
		03932 => "11111111",
		03933 => "11111111",
		03934 => "11111111",
		03935 => "11111111",
		03936 => "11111111",
		03937 => "11111111",
		03938 => "11111111",
		03939 => "11111111",
		03940 => "11111111",
		03941 => "11111111",
		03942 => "11111111",
		03943 => "11111111",
		03944 => "11111111",
		03945 => "11111111",
		03946 => "11111111",
		03947 => "11111111",
		03948 => "11111111",
		03949 => "11111111",
		03950 => "11111111",
		03951 => "11111111",
		03952 => "11111111",
		03953 => "11111111",
		03954 => "11111111",
		03955 => "11111111",
		03956 => "11111111",
		03957 => "11111111",
		03958 => "11111111",
		03959 => "11111111",
		03960 => "11111111",
		03961 => "11111111",
		03962 => "11111111",
		03963 => "11111111",
		03964 => "11111111",
		03965 => "11111111",
		03966 => "11111111",
		03967 => "11111111",
		03968 => "11111111",
		03969 => "11111111",
		03970 => "11111111",
		03971 => "11111111",
		03972 => "11111111",
		03973 => "11111111",
		03974 => "11111111",
		03975 => "11111111",
		03976 => "11111111",
		03977 => "11111111",
		03978 => "11111111",
		03979 => "11111111",
		03980 => "11111111",
		03981 => "11111111",
		03982 => "11111111",
		03983 => "11111111",
		03984 => "11111111",
		03985 => "11111111",
		03986 => "11111111",
		03987 => "11111111",
		03988 => "11111111",
		03989 => "11111111",
		03990 => "11111111",
		03991 => "11111111",
		03992 => "11111111",
		03993 => "11111111",
		03994 => "11111111",
		03995 => "11111111",
		03996 => "11111111",
		03997 => "11111111",
		03998 => "11111111",
		03999 => "11111111",
		04000 => "11111111",
		04001 => "11111111",
		04002 => "11111111",
		04003 => "11111111",
		04004 => "11111111",
		04005 => "11111111",
		04006 => "11111111",
		04007 => "11111111",
		04008 => "11111111",
		04009 => "11111111",
		04010 => "11111111",
		04011 => "11111111",
		04012 => "11111111",
		04013 => "11111111",
		04014 => "11111111",
		04015 => "11111111",
		04016 => "11111111",
		04017 => "11111111",
		04018 => "11111111",
		04019 => "11111111",
		04020 => "11111111",
		04021 => "11111111",
		04022 => "11111111",
		04023 => "11111111",
		04024 => "11111111",
		04025 => "11111111",
		04026 => "11111111",
		04027 => "11111111",
		04028 => "11111111",
		04029 => "11111111",
		04030 => "11111111",
		04031 => "11111111",
		04032 => "11111111",
		04033 => "11111111",
		04034 => "11111111",
		04035 => "11111111",
		04036 => "11111111",
		04037 => "11111111",
		04038 => "11111111",
		04039 => "11111111",
		04040 => "11111111",
		04041 => "11111111",
		04042 => "11111111",
		04043 => "11111111",
		04044 => "11111111",
		04045 => "11111111",
		04046 => "11111111",
		04047 => "11111111",
		04048 => "11111111",
		04049 => "11111111",
		04050 => "11111111",
		04051 => "11111111",
		04052 => "11111111",
		04053 => "11111111",
		04054 => "11111111",
		04055 => "11111111",
		04056 => "11111111",
		04057 => "11111111",
		04058 => "11111111",
		04059 => "11111111",
		04060 => "11111111",
		04061 => "11111111",
		04062 => "11111111",
		04063 => "11111111",
		04064 => "11111111",
		04065 => "11111111",
		04066 => "11111111",
		04067 => "11111111",
		04068 => "11111111",
		04069 => "11111111",
		04070 => "11111111",
		04071 => "11111111",
		04072 => "11111111",
		04073 => "11111111",
		04074 => "11111111",
		04075 => "11111111",
		04076 => "11111111",
		04077 => "11111111",
		04078 => "11111111",
		04079 => "11111111",
		04080 => "11111111",
		04081 => "11111111",
		04082 => "11111111",
		04083 => "11111111",
		04084 => "11111111",
		04085 => "11111111",
		04086 => "11111111",
		04087 => "11111111",
		04088 => "11111111",
		04089 => "11111111",
		04090 => "11111111",
		04091 => "11111111",
		04092 => "11111111",
		04093 => "11111111",
		04094 => "11111111",
		04095 => "11111111",
		OTHERS=> "11111111"
		);

BEGIN
  A <= (                        A11 & A10 & A09 & A08 &
        A07 & A06 & A05 & A04 & A03 & A02 & A01 & A00 );
  --
  PROCESS( CS, A )
  BEGIN
    if (CS = '1') then
          D <= ROM_Cells(to_integer(unsigned(A))); -- READ condition
    else  D <= (others => '0');                    -- Chip Select Off
    end if;
  END PROCESS;
  --
  D07 <= D(7); D06 <= D(6); D05 <= D(5); D04 <= D(4);
  D03 <= D(3); D02 <= D(2); D01 <= D(1); D00 <= D(0);
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY NOT_gate IS
  PORT( I: IN std_logic;
  	O: OUT std_logic );
END NOT_gate;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF NOT_gate IS
BEGIN
  O <= (not I);
END behavioral;



--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY AND2_gate IS
  PORT( I0,I1: IN std_logic;
        O: OUT std_logic );
END AND2_gate;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF AND2_gate IS
BEGIN
  O <= (I0 and I1);
END behavioral;


--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY Multiplexer_2_1 IS

  PORT( I0: IN  std_logic;
        I1: IN  std_logic;
        S0: IN  std_logic;
         Q: OUT std_logic );
END Multiplexer_2_1;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF Multiplexer_2_1 IS
BEGIN
  Q <= I0 when (S0 = '0') else
       I1 when (S0 = '1') else 'X';
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY BusMultiplexer21_8 IS

  PORT( Q_07: OUT std_logic;
        Q_06: OUT std_logic;
        Q_05: OUT std_logic;
        Q_04: OUT std_logic;
        Q_03: OUT std_logic;
        Q_02: OUT std_logic;
        Q_01: OUT std_logic;
        Q_00: OUT std_logic;
        I0_07: IN  std_logic;
        I0_06: IN  std_logic;
        I0_05: IN  std_logic;
        I0_04: IN  std_logic;
        I0_03: IN  std_logic;
        I0_02: IN  std_logic;
        I0_01: IN  std_logic;
        I0_00: IN  std_logic;
        I1_07: IN  std_logic;
        I1_06: IN  std_logic;
        I1_05: IN  std_logic;
        I1_04: IN  std_logic;
        I1_03: IN  std_logic;
        I1_02: IN  std_logic;
        I1_01: IN  std_logic;
        I1_00: IN  std_logic;
        S0  :  IN  std_logic );
END BusMultiplexer21_8;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF BusMultiplexer21_8 IS
BEGIN
  Q_07 <= I0_07 when (S0 = '0') else
          I1_07 when (S0 = '1') else 'X';
  Q_06 <= I0_06 when (S0 = '0') else
          I1_06 when (S0 = '1') else 'X';
  Q_05 <= I0_05 when (S0 = '0') else
          I1_05 when (S0 = '1') else 'X';
  Q_04 <= I0_04 when (S0 = '0') else
          I1_04 when (S0 = '1') else 'X';
  Q_03 <= I0_03 when (S0 = '0') else
          I1_03 when (S0 = '1') else 'X';
  Q_02 <= I0_02 when (S0 = '0') else
          I1_02 when (S0 = '1') else 'X';
  Q_01 <= I0_01 when (S0 = '0') else
          I1_01 when (S0 = '1') else 'X';
  Q_00 <= I0_00 when (S0 = '0') else
          I1_00 when (S0 = '1') else 'X';
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY BusMultiplexer21_16 IS

  PORT( Q_15: OUT std_logic;
        Q_14: OUT std_logic;
        Q_13: OUT std_logic;
        Q_12: OUT std_logic;
        Q_11: OUT std_logic;
        Q_10: OUT std_logic;
        Q_09: OUT std_logic;
        Q_08: OUT std_logic;
        Q_07: OUT std_logic;
        Q_06: OUT std_logic;
        Q_05: OUT std_logic;
        Q_04: OUT std_logic;
        Q_03: OUT std_logic;
        Q_02: OUT std_logic;
        Q_01: OUT std_logic;
        Q_00: OUT std_logic;
        I0_15: IN  std_logic;
        I0_14: IN  std_logic;
        I0_13: IN  std_logic;
        I0_12: IN  std_logic;
        I0_11: IN  std_logic;
        I0_10: IN  std_logic;
        I0_09: IN  std_logic;
        I0_08: IN  std_logic;
        I0_07: IN  std_logic;
        I0_06: IN  std_logic;
        I0_05: IN  std_logic;
        I0_04: IN  std_logic;
        I0_03: IN  std_logic;
        I0_02: IN  std_logic;
        I0_01: IN  std_logic;
        I0_00: IN  std_logic;
        I1_15: IN  std_logic;
        I1_14: IN  std_logic;
        I1_13: IN  std_logic;
        I1_12: IN  std_logic;
        I1_11: IN  std_logic;
        I1_10: IN  std_logic;
        I1_09: IN  std_logic;
        I1_08: IN  std_logic;
        I1_07: IN  std_logic;
        I1_06: IN  std_logic;
        I1_05: IN  std_logic;
        I1_04: IN  std_logic;
        I1_03: IN  std_logic;
        I1_02: IN  std_logic;
        I1_01: IN  std_logic;
        I1_00: IN  std_logic;
        S0  :  IN  std_logic );
END BusMultiplexer21_16;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF BusMultiplexer21_16 IS
BEGIN
  Q_15 <= I0_15 when (S0 = '0') else
          I1_15 when (S0 = '1') else 'X';
  Q_14 <= I0_14 when (S0 = '0') else
          I1_14 when (S0 = '1') else 'X';
  Q_13 <= I0_13 when (S0 = '0') else
          I1_13 when (S0 = '1') else 'X';
  Q_12 <= I0_12 when (S0 = '0') else
          I1_12 when (S0 = '1') else 'X';
  Q_11 <= I0_11 when (S0 = '0') else
          I1_11 when (S0 = '1') else 'X';
  Q_10 <= I0_10 when (S0 = '0') else
          I1_10 when (S0 = '1') else 'X';
  Q_09 <= I0_09 when (S0 = '0') else
          I1_09 when (S0 = '1') else 'X';
  Q_08 <= I0_08 when (S0 = '0') else
          I1_08 when (S0 = '1') else 'X';
  Q_07 <= I0_07 when (S0 = '0') else
          I1_07 when (S0 = '1') else 'X';
  Q_06 <= I0_06 when (S0 = '0') else
          I1_06 when (S0 = '1') else 'X';
  Q_05 <= I0_05 when (S0 = '0') else
          I1_05 when (S0 = '1') else 'X';
  Q_04 <= I0_04 when (S0 = '0') else
          I1_04 when (S0 = '1') else 'X';
  Q_03 <= I0_03 when (S0 = '0') else
          I1_03 when (S0 = '1') else 'X';
  Q_02 <= I0_02 when (S0 = '0') else
          I1_02 when (S0 = '1') else 'X';
  Q_01 <= I0_01 when (S0 = '0') else
          I1_01 when (S0 = '1') else 'X';
  Q_00 <= I0_00 when (S0 = '0') else
          I1_00 when (S0 = '1') else 'X';
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Adder_16 IS

  PORT( CIN: IN  std_logic;
        COUT:OUT std_logic;
        OVF: OUT std_logic;
        A15: IN  std_logic;
        A14: IN  std_logic;
        A13: IN  std_logic;
        A12: IN  std_logic;
        A11: IN  std_logic;
        A10: IN  std_logic;
        A9:  IN  std_logic;
        A8:  IN  std_logic;
        A7:  IN  std_logic;
        A6:  IN  std_logic;
        A5:  IN  std_logic;
        A4:  IN  std_logic;
        A3:  IN  std_logic;
        A2:  IN  std_logic;
        A1:  IN  std_logic;
        A0:  IN  std_logic;
        B15: IN  std_logic;
        B14: IN  std_logic;
        B13: IN  std_logic;
        B12: IN  std_logic;
        B11: IN  std_logic;
        B10: IN  std_logic;
        B9:  IN  std_logic;
        B8:  IN  std_logic;
        B7:  IN  std_logic;
        B6:  IN  std_logic;
        B5:  IN  std_logic;
        B4:  IN  std_logic;
        B3:  IN  std_logic;
        B2:  IN  std_logic;
        B1:  IN  std_logic;
        B0:  IN  std_logic;
        F15: OUT std_logic;
        F14: OUT std_logic;
        F13: OUT std_logic;
        F12: OUT std_logic;
        F11: OUT std_logic;
        F10: OUT std_logic;
        F9:  OUT std_logic;
        F8:  OUT std_logic;
        F7:  OUT std_logic;
        F6:  OUT std_logic;
        F5:  OUT std_logic;
        F4:  OUT std_logic;
        F3:  OUT std_logic;
        F2:  OUT std_logic;
        F1:  OUT std_logic;
        F0:  OUT std_logic );
END Adder_16;
--------------------------------------------------------------------
ARCHITECTURE behavioral OF Adder_16 IS
BEGIN
  Add16: PROCESS( A15, A14, A13, A12, A11, A10, A9, A8,
                  A7,  A6,  A5,  A4,  A3,  A2,  A1, A0,
                  B15, B14, B13, B12, B11, B10, B9, B8,
                  B7,  B6,  B5,  B4,  B3,  B2,  B1, B0,
                  CIN )
  variable A : unsigned(16 downto 0 );
  variable B : unsigned(16 downto 0 );
  variable Ar: unsigned(16 downto 0 );  --(without the sign bit)
  variable Br: unsigned(16 downto 0 );
  variable F : unsigned(16 downto 0 );
  BEGIN
    A := ('0'& A15 & A14 & A13 & A12 & A11 & A10 & A9 & A8
             & A7  & A6  & A5  & A4  & A3  & A2  & A1 & A0);
    B := ('0'& B15 & B14 & B13 & B12 & B11 & B10 & B9 & B8
             & B7  & B6  & B5  & B4  & B3  & B2  & B1 & B0);
    --
    Ar:= ('0'&'0' & A14 & A13 & A12 & A11 & A10 & A9 & A8  --(without the sign bit)
             & A7 & A6  & A5  & A4  & A3  & A2  & A1 & A0);
    Br:= ('0'&'0' & B14 & B13 & B12 & B11 & B10 & B9 & B8
             & B7 & B6  & B5  & B4  & B3  & B2  & B1 & B0);
    --
    if    (CIN = '0') then  F := Ar + Br;
    elsif (CIN = '1') then  F := Ar + Br + 1;
    else                    F := (others =>'X');  -- (CIN: Unknown)
    END IF;
    --
    OVF  <= ((not F(15)) and (    A(15)) and (    B(15))) or
            ((    F(15)) and (not A(15)) and (not B(15)));
    COUT <= (A(15) and B(15)) or
            (A(15) and F(15)) or
            (B(15) and F(15));
    F15  <= (A(15) xor B(15)) xor F(15);
    F14  <=  F(14);
    F13  <=  F(13);
    F12  <=  F(12);
    F11  <=  F(11);
    F10  <=  F(10);
    F9   <=  F(9);
    F8   <=  F(8);
    F7   <=  F(7);
    F6   <=  F(6);
    F5   <=  F(5);
    F4   <=  F(4);
    F3   <=  F(3);
    F2   <=  F(2);
    F1   <=  F(1);
    F0   <=  F(0);
  END PROCESS;
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Multiplier_8x8 IS

  PORT( SNA:  IN  std_logic;
        SNB:  IN  std_logic;
        A07:  IN  std_logic;
        A06:  IN  std_logic;
        A05:  IN  std_logic;
        A04:  IN  std_logic;
        A03:  IN  std_logic;
        A02:  IN  std_logic;
        A01:  IN  std_logic;
        A00:  IN  std_logic;
        B07:  IN  std_logic;
        B06:  IN  std_logic;
        B05:  IN  std_logic;
        B04:  IN  std_logic;
        B03:  IN  std_logic;
        B02:  IN  std_logic;
        B01:  IN  std_logic;
        B00:  IN  std_logic;
		  M15:  OUT std_logic;
		  M14:  OUT std_logic;
		  M13:  OUT std_logic;
		  M12:  OUT std_logic;
		  M11:  OUT std_logic;
		  M10:  OUT std_logic;
		  M09:  OUT std_logic;
		  M08:  OUT std_logic;
		  M07:  OUT std_logic;
        M06:  OUT std_logic;
        M05:  OUT std_logic;
        M04:  OUT std_logic;
        M03:  OUT std_logic;
        M02:  OUT std_logic;
        M01:  OUT std_logic;
        M00:  OUT std_logic );
END Multiplier_8x8;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF Multiplier_8x8 IS

	signal sign: std_logic;
	signal A_in: STD_LOGIC_VECTOR ( 7 downto 0 ); 
	signal B_in: STD_LOGIC_VECTOR ( 7 downto 0 ); 
	signal AM  : STD_LOGIC_VECTOR ( 7 downto 0 ); 
	signal BM  : STD_LOGIC_VECTOR ( 7 downto 0 ); 
	signal R   : STD_LOGIC_VECTOR (15 downto 0 );
	
BEGIN
   A_in <= ( A07 & A06 & A05 & A04 & A03 & A02 & A01 & A00 );
	B_in <= ( B07 & B06 & B05 & B04 & B03 & B02 & B01 & B00 );

   AM <= A_in 	when (SNA = '0') or (A07 = '0') 
					else std_logic_vector( unsigned(not(A_in))+1 );
	BM <= B_in	when (SNB = '0') or (B07 = '0') 
					else std_logic_vector( unsigned(not(B_in))+1 );

	sign <=	(A07 and SNA) xor (B07 and SNB);  -- sign of result
	R <= 	std_logic_vector( unsigned(AM) * unsigned(BM) ) when sign = '0' 
			else std_logic_vector( not(unsigned(AM) * unsigned(BM)) +1);
	
	M15 <= R(15);	M14 <= R(14);	M13 <= R(13);	M12 <= R(12);	
	M11 <= R(11);	M10 <= R(10);	M09 <= R(09);	M08 <= R(08);
	M07 <= R(7);	M06 <= R(6);	M05 <= R(5);	M04 <= R(4);
	M03 <= R(3);	M02 <= R(2);	M01 <= R(1);	M00 <= R(0);
	
END behavioral;
--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY DpetFF IS
  PORT(  D, Ck   : IN std_logic;
         nCL, nPR: IN std_logic;
         Q, nQ   : OUT std_logic );
END DpetFF;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF DpetFF IS 
BEGIN
  Dff: PROCESS( Ck, nCL, nPR ) 
  BEGIN
    if    (nCL = '0') and (nPR = '0') then  Q <= 'X';  nQ <= 'X';
    elsif (nCL = '0') and (nPR = '1') then  Q <= '0';  nQ <= '1';
    elsif (nCL = '1') and (nPR = '0') then  Q <= '1';  nQ <= '0';
    elsif (nCL = '1') and (nPR = '1') then
      if (Ck'event) AND (Ck='1') THEN -- Positive Edge -----------
                                            Q <=  D;   nQ <= not D;
      END IF;
    else                                    Q <= 'X';  nQ <= 'X';
    END IF;
  END PROCESS; 
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY EpetFF IS
  PORT(  D, E, Ck: IN std_logic;
         nCL, nPR: IN std_logic;
         Q, nQ   : OUT std_logic );
END EpetFF;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF EpetFF IS 
BEGIN
  Eff: PROCESS( Ck, nCL, nPR )
  BEGIN
    if    (nCL = '0') and (nPR = '0') then  Q <= 'X';  nQ <= 'X';
    elsif (nCL = '0') and (nPR = '1') then  Q <= '0';  nQ <= '1';
    elsif (nCL = '1') and (nPR = '0') then  Q <= '1';  nQ <= '0';
    elsif (nCL = '1') and (nPR = '1') then
      if (Ck'event) AND (Ck='1') THEN -- Positive Edge -----------
        if (E = '1') then                   Q <=  D;   nQ <= not D;
        elsif not(E = '0') then             Q <= 'X';  nQ <= 'X';
        END IF;
      END IF;
    else                                    Q <= 'X';  nQ <= 'X';
    END IF;
  END PROCESS;
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Counter8b IS
  PORT( Ck : IN std_logic;
        nCL: IN std_logic;
        LD : IN std_logic;
        ENP: IN std_logic;
        ENT: IN std_logic;
        UD : IN std_logic;

        P7 : IN std_logic;
        P6 : IN std_logic;
        P5 : IN std_logic;
        P4 : IN std_logic;
        P3 : IN std_logic;
        P2 : IN std_logic;
        P1 : IN std_logic;
        P0 : IN std_logic;

        Q7 : OUT std_logic;
        Q6 : OUT std_logic;
        Q5 : OUT std_logic;
        Q4 : OUT std_logic;
        Q3 : OUT std_logic;
        Q2 : OUT std_logic;
        Q1 : OUT std_logic;
        Q0 : OUT std_logic;

        Tc : OUT std_logic );
END Counter8b;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF Counter8b IS
BEGIN
  Count8b: PROCESS( Ck, nCL, ENP, ENT, UD )
  variable aCnt: unsigned( 7 downto 0 );
  BEGIN
    if    (nCL = '0') then                aCnt := (others =>'0');
    elsif (nCL = '1') then
      if (Ck'event) AND (Ck='1') then
        if    (LD = '1') then             aCnt := (P7 & P6 & P5 & P4 & P3 & P2 & P1 & P0); -- Load
        elsif (LD = '0') then
          if  (ENP = '1') and (ENT = '1')then
            if    (UD = '1') then
              if (aCnt < "11111111") then aCnt := aCnt + 1;
              else                        aCnt := (others =>'0');
              end if;
            elsif (UD = '0') then
              if (aCnt > "00000000") then aCnt := aCnt - 1;
              else                        aCnt := (others =>'1');
              end if;
            else                          aCnt := (others =>'X'); -- (UD: Unknown)
            END IF;
          elsif not((ENP ='0')or
                    (ENT ='0') ) then     aCnt := (others =>'X'); -- (EN: Unknown)
          END IF;
        else                              aCnt := (others =>'X'); -- (LD: Unknown)
        END IF;
      END IF;
    else                                  aCnt := (others =>'X'); -- (nCL: Unknown)
    END IF;
    --
    Tc <= ENT and (    (aCnt(7) and aCnt(6) and aCnt(5) and aCnt(4) and aCnt(3) and aCnt(2) and aCnt(1) and aCnt(0) and UD) or
                   (not(aCnt(7) or  aCnt(6) or  aCnt(5) or  aCnt(4) or  aCnt(3) or  aCnt(2) or  aCnt(1) or  aCnt(0) or  UD))  );
    --
    Q7 <= aCnt(7);
    Q6 <= aCnt(6);
    Q5 <= aCnt(5);
    Q4 <= aCnt(4);
    Q3 <= aCnt(3);
    Q2 <= aCnt(2);
    Q1 <= aCnt(1);
    Q0 <= aCnt(0);
    --
  END PROCESS;
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Counter16 IS
  PORT( Ck : IN std_logic;
        nCL: IN std_logic;
        LD : IN std_logic;
        ENP: IN std_logic;
        ENT: IN std_logic;
        UD : IN std_logic;

        P15: IN std_logic;
        P14: IN std_logic;
        P13: IN std_logic;
        P12: IN std_logic;
        P11: IN std_logic;
        P10: IN std_logic;
        P9 : IN std_logic;
        P8 : IN std_logic;

        P7 : IN std_logic;
        P6 : IN std_logic;
        P5 : IN std_logic;
        P4 : IN std_logic;
        P3 : IN std_logic;
        P2 : IN std_logic;
        P1 : IN std_logic;
        P0 : IN std_logic;

        Q15: OUT std_logic;
        Q14: OUT std_logic;
        Q13: OUT std_logic;
        Q12: OUT std_logic;
        Q11: OUT std_logic;
        Q10: OUT std_logic;
        Q9 : OUT std_logic;
        Q8 : OUT std_logic;

        Q7 : OUT std_logic;
        Q6 : OUT std_logic;
        Q5 : OUT std_logic;
        Q4 : OUT std_logic;
        Q3 : OUT std_logic;
        Q2 : OUT std_logic;
        Q1 : OUT std_logic;
        Q0 : OUT std_logic;

        Tc : OUT std_logic );
END Counter16;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF Counter16 IS
BEGIN
  Count16: PROCESS( Ck, nCL, ENP, ENT, UD )
  variable aCnt: unsigned( 15 downto 0 );
  BEGIN
    if    (nCL = '0') then                        aCnt := (others =>'0');
    elsif (nCL = '1') then
      if (Ck'event) AND (Ck='1') then
        if    (LD = '1') then                     aCnt := (P15 & P14 & P13 & P12 & P11 & P10 & P9 & P8 &  -- Load
                                                           P7  & P6  & P5  & P4  & P3  & P2  & P1 & P0);
        elsif (LD = '0') then
          if  (ENP = '1') and (ENT = '1')then
            if    (UD = '1') then
              if (aCnt < "1111111111111111") then aCnt := aCnt + 1;
              else                                aCnt := (others =>'0');
              end if;
            elsif (UD = '0') then
              if (aCnt > "0000000000000000") then aCnt := aCnt - 1;
              else                                aCnt := (others =>'1');
              end if;
            else                                  aCnt := (others =>'X'); -- (UD: Unknown)
            END IF;
          elsif not((ENP ='0')or
                    (ENT ='0') ) then             aCnt := (others =>'X'); -- (EN: Unknown)
          END IF;
        else                                      aCnt := (others =>'X'); -- (LD: Unknown)
        END IF;
      END IF;
    else                                          aCnt := (others =>'X'); -- (nCL: Unknown)
    END IF;
    --
    Tc <= ENT and (   (aCnt(15) and aCnt(14) and aCnt(13) and aCnt(12) and aCnt(11) and aCnt(10) and aCnt(9) and aCnt(8) and
                       aCnt( 7) and aCnt( 6) and aCnt( 5) and aCnt( 4) and aCnt( 3) and aCnt( 2) and aCnt(1) and aCnt(0) and UD) or
                  (not(aCnt(15) or  aCnt(14) or  aCnt(13) or  aCnt(12) or  aCnt(11) or  aCnt(10) or  aCnt(9) or  aCnt(8) or
                       aCnt( 7) or  aCnt( 6) or  aCnt( 5) or  aCnt( 4) or  aCnt( 3) or  aCnt( 2) or  aCnt(1) or  aCnt(0) or UD))   );
    --
    Q15 <= aCnt(15);
    Q14 <= aCnt(14);
    Q13 <= aCnt(13);
    Q12 <= aCnt(12);
    Q11 <= aCnt(11);
    Q10 <= aCnt(10);
    Q9  <= aCnt(9);
    Q8  <= aCnt(8);
    Q7  <= aCnt(7);
    Q6  <= aCnt(6);
    Q5  <= aCnt(5);
    Q4  <= aCnt(4);
    Q3  <= aCnt(3);
    Q2  <= aCnt(2);
    Q1  <= aCnt(1);
    Q0  <= aCnt(0);
    --
  END PROCESS;
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY PiPoE8b IS
  PORT( Ck : IN std_logic;
        nCL: IN std_logic;
        E  : IN std_logic;
        P7 : IN std_logic;
        P6 : IN std_logic;
        P5 : IN std_logic;
        P4 : IN std_logic;
        P3 : IN std_logic;
        P2 : IN std_logic;
        P1 : IN std_logic;
        P0 : IN std_logic;
        Q7 : OUT std_logic;
        Q6 : OUT std_logic;
        Q5 : OUT std_logic;
        Q4 : OUT std_logic;
        Q3 : OUT std_logic;
        Q2 : OUT std_logic;
        Q1 : OUT std_logic;
        Q0 : OUT std_logic );
END PiPoE8b;


--------------------------------------------------------------------
ARCHITECTURE behavioral OF PiPoE8b IS
BEGIN
  RegPiPoE8b: PROCESS( Ck, nCL )
    variable aReg: std_logic_vector( 7 downto 0 );
  BEGIN
    if    (nCL = '0') then    aReg := (others =>'0');
    elsif (nCL = '1') then
      if (Ck'event) AND (Ck='1') THEN -- Positive Edge -----------
        if (E = '1') then
                aReg := (P7 & P6 & P5 & P4 & P3 & P2 & P1 & P0);
        elsif not(E = '0') then
                aReg := (others =>'X');
        END IF;
      END IF;
    else        aReg := (others =>'X');
    END IF;

    Q7 <= aReg(7);
    Q6 <= aReg(6);
    Q5 <= aReg(5);
    Q4 <= aReg(4);
    Q3 <= aReg(3);
    Q2 <= aReg(2);
    Q1 <= aReg(1);
    Q0 <= aReg(0);

  END PROCESS;
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY PiPoE16 IS
  PORT( Ck : IN std_logic;
        nCL: IN std_logic;
        E  : IN std_logic;
        P15: IN std_logic;
        P14: IN std_logic;
        P13: IN std_logic;
        P12: IN std_logic;
        P11: IN std_logic;
        P10: IN std_logic;
        P9 : IN std_logic;
        P8 : IN std_logic;
        P7 : IN std_logic;
        P6 : IN std_logic;
        P5 : IN std_logic;
        P4 : IN std_logic;
        P3 : IN std_logic;
        P2 : IN std_logic;
        P1 : IN std_logic;
        P0 : IN std_logic;
        Q15: OUT std_logic;
        Q14: OUT std_logic;
        Q13: OUT std_logic;
        Q12: OUT std_logic;
        Q11: OUT std_logic;
        Q10: OUT std_logic;
        Q9 : OUT std_logic;
        Q8 : OUT std_logic;
        Q7 : OUT std_logic;
        Q6 : OUT std_logic;
        Q5 : OUT std_logic;
        Q4 : OUT std_logic;
        Q3 : OUT std_logic;
        Q2 : OUT std_logic;
        Q1 : OUT std_logic;
        Q0 : OUT std_logic );
END PiPoE16;


--------------------------------------------------------------------
ARCHITECTURE behavioral OF PiPoE16 IS
BEGIN
  RegPiPoE16: PROCESS( Ck, nCL )
    variable aReg: std_logic_vector( 15 downto 0 );
  BEGIN
    if    (nCL = '0') then    aReg := (others =>'0');
    elsif (nCL = '1') then
      if (Ck'event) AND (Ck='1') THEN -- Positive Edge -----------
        if (E = '1') then
                aReg := (P15 & P14 & P13 & P12 & P11 & P10 & P9 & P8 &
                         P7  & P6  & P5  & P4  & P3  & P2  & P1 & P0);
        elsif not(E = '0') then
                aReg := (others =>'X');
        END IF;
      END IF;
    else        aReg := (others =>'X');
    END IF;

    Q15 <= aReg(15);
    Q14 <= aReg(14);
    Q13 <= aReg(13);
    Q12 <= aReg(12);
    Q11 <= aReg(11);
    Q10 <= aReg(10);
    Q9  <= aReg(9);
    Q8  <= aReg(8);
    Q7  <= aReg(7);
    Q6  <= aReg(6);
    Q5  <= aReg(5);
    Q4  <= aReg(4);
    Q3  <= aReg(3);
    Q2  <= aReg(2);
    Q1  <= aReg(1);
    Q0  <= aReg(0);

  END PROCESS;
END behavioral;

--------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

ENTITY PiSoE16 IS
  PORT( Ck : IN std_logic;
        nCL: IN std_logic;
        E  : IN std_logic;
        LD : IN std_logic;
        P15: IN std_logic;
        P14: IN std_logic;
        P13: IN std_logic;
        P12: IN std_logic;
        P11: IN std_logic;
        P10: IN std_logic;
        P9 : IN std_logic;
        P8 : IN std_logic;
        P7 : IN std_logic;
        P6 : IN std_logic;
        P5 : IN std_logic;
        P4 : IN std_logic;
        P3 : IN std_logic;
        P2 : IN std_logic;
        P1 : IN std_logic;
        P0 : IN std_logic;
        Q0 : OUT std_logic );
END PiSoE16;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF PiSoE16 IS
BEGIN
  RegPiSoE16: PROCESS( Ck, nCL, LD )
  variable aReg: std_logic_vector(15 downto 0 );
  BEGIN
    if    (nCL = '0') then    aReg := (others =>'0');
    elsif (nCL = '1') then
      if (Ck'event) AND (Ck='1') THEN -- Positive Edge -----------
        if  (LD = '1') then
                  aReg := (P15 & P14 & P13 & P12 & P11 & P10 & P9 & P8 &
                           P7  & P6  & P5  & P4  & P3  & P2  & P1 & P0);
        elsif(LD = '0') then
          if (E = '1') then
                  aReg := ('0'     & aReg(15) & aReg(14) & aReg(13) & aReg(12) & aReg(11) & aReg(10) & aReg(9) &
                           aReg(8) & aReg(7)  & aReg(6)  & aReg(5)  & aReg(4)  & aReg(3)  & aReg(2)  & aReg(1));
          elsif not(E = '0') then
                  aReg := (others =>'X');
          END IF;
        else      aReg := (others =>'X');
        END IF;
      END IF;
    else          aReg := (others =>'X');
    END IF;
    ----------------
    Q0 <= aReg(0);
  END PROCESS;
END behavioral;

--------------------------------------------------------------------
LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY SSRAM256x8 IS           -- Synchronous Static RAM 256 x 8
  PORT( CK  : IN  std_logic;
        CS  : IN  std_logic;
        WE  : IN  std_logic;
        A00 : IN  std_logic;   -- ADR 14..0 (32K)
        A01 : IN  std_logic;
        A02 : IN  std_logic;
        A03 : IN  std_logic;
        A04 : IN  std_logic;
        A05 : IN  std_logic;
        A06 : IN  std_logic;
        A07 : IN  std_logic;
        D00 : IN  std_logic;   -- Data Input 07..00 (8-bits)
        D01 : IN  std_logic;
        D02 : IN  std_logic;
        D03 : IN  std_logic;
        D04 : IN  std_logic;
        D05 : IN  std_logic;
        D06 : IN  std_logic;
        D07 : IN  std_logic;
        Q00 : OUT std_logic;   -- Data Output 07..00 (8-bits)
        Q01 : OUT std_logic;
        Q02 : OUT std_logic;
        Q03 : OUT std_logic;
        Q04 : OUT std_logic;
        Q05 : OUT std_logic;
        Q06 : OUT std_logic;
        Q07 : OUT std_logic );
END SSRAM256x8;

--------------------------------------------------------------------
ARCHITECTURE behavioral OF SSRAM256x8 IS
  --
  type RAM_Array is array (0 to 255) of std_logic_vector(7 downto 0);
  --
  SIGNAL RAM_Cells: RAM_Array;
  SIGNAL A : std_logic_vector( 7 downto 0);
  SIGNAL AR: std_logic_vector( 7 downto 0);
  SIGNAL Q : std_logic_vector( 7 downto 0);

BEGIN
  A <= (A07 & A06 & A05 & A04 & A03 & A02 & A01 & A00);
  --
  PROCESS( CK )
  BEGIN
    if (CS = '1') then
      if (CK'event and (CK = '1')) then
        if (WE = '1') then
             RAM_Cells(to_integer(unsigned(A))) <=( D07 & D06 & D05 & D04 &
                                                    D03 & D02 & D01 & D00 );
        end if;
        AR <= A;
      end if;
    end if;
  END PROCESS;
  --
  Q <= RAM_Cells(to_integer(unsigned(AR))) when (CS = '1') else
       (others => '0');
  Q07 <= Q(7); Q06 <= Q(6); Q05 <= Q(5); Q04 <= Q(4);
  Q03 <= Q(3); Q02 <= Q(2); Q01 <= Q(1); Q00 <= Q(0);
END behavioral;


